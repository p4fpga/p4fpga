method forward_table_add_entry=ingress.forward_table_add_entry;
