method forward_table_add_entry = prog.forward_table_add_entry;
