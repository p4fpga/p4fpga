
typedef enum {
  NOP,
  FORWARD
} RouteActionT deriving (Bits, Eq);


