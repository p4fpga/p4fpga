import Ethernet::*;
