method forward_add_entry = prog.forward_add_entry;
method ipv4_lpm_add_entry = prog.ipv4_lpm_add_entry;
method t_opti_update_add_entry = prog.t_opti_update_add_entry;
method t_reply_client_add_entry = prog.t_reply_client_add_entry;
method t_req_fix_add_entry = prog.t_req_fix_add_entry;
method t_req_pass1_add_entry = prog.t_req_pass1_add_entry;
method t_store_update_add_entry = prog.t_store_update_add_entry;
method send_frame_add_entry = prog.send_frame_add_entry;
