
typedef enum {
  NOP,
  FORWARD
} FwdTblActionT deriving (Bits, Eq);


