method forward_table_add_entry = prog.forward_table_add_entry;
method table_1_add_entry = prog.table_1_add_entry;
method table_2_add_entry = prog.table_2_add_entry;
method table_3_add_entry = prog.table_3_add_entry;
method table_4_add_entry = prog.table_4_add_entry;
method table_5_add_entry = prog.table_5_add_entry;
method table_6_add_entry = prog.table_6_add_entry;
method table_7_add_entry = prog.table_7_add_entry;
