method Action forward_table_add_entry(ForwardTableReqT key, ForwardTableRspT val);
method Action test_tbl_add_entry(TestTblReqT key, TestTblRspT val);
