
Reg#(Bit#(32)) test <- mkReg(0);
