method forward_add_entry = prog.forward_add_entry;
method ipv4_lpm_add_entry = prog.ipv4_lpm_add_entry;
method send_frame_add_entry = prog.send_frame_add_entry;
