import Library::*;

export Ingress(..), mkIngress;
export Egress(..), mkEgress;

`include "ControlGenerated.bsv"
