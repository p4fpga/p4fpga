method Action forward_table_add_entry(ForwardTableReqT key, ForwardTableRspT val);
