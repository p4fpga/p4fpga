import StructGenerated::*;
