method Action forward_add_entry(ForwardReqT key, ForwardRspT nhop_ipv4);
