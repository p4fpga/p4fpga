method Action forward_add_entry(ForwardReqSize key, ForwardRspSize value);
method Action ipv4_lpm_add_entry(Ipv4LpmReqSize key, Ipv4LpmRspSize value);
method Action send_frame_add_entry(SendFrameReqSize key, SendFrameRspSize value);
