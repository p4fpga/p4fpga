
typedef enum {
  NOP,
  FORWARD
} RoutingActionT deriving (Bits, Eq);


