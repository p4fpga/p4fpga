import Ethernet::*;
typedef union tagged {
  struct {
    PacketInstance pkt;
  } DropReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) stats_metadata$flow_map_index;
  } GetSenderIpReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(2) stats_metadata$flow_map_index;
  } IncreaseMincwndReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) stats_metadata$flow_map_index;
  } LookupFlowMapReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) stats_metadata$flow_map_index;
  } LookupFlowMapReverseReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) options_wscale$wscale;
    Bit#(2) stats_metadata$flow_map_index;
    Bit#(16) options_mss$mss;
    Bit#(32) ipv4$dstAddr;
  } RecordIpReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) runtime_smac_48;
  } RewriteMacReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) stats_metadata$flow_map_index;
    Bit#(32) tcp$seqNo;
    Bit#(48) intrinsic_metadata$ingress_global_timestamp;
  } SampleNewRttReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) stats_metadata$flow_map_index;
    Bit#(32) stats_metadata$senderIP;
    Bit#(32) ipv4$srcAddr;
    Bit#(32) ipv4$dstAddr;
  } SaveSourceIpReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) runtime_dmac_48;
  } SetDmacReqT;
  struct {
    PacketInstance pkt;
    Bit#(9) runtime_port_9;
    Bit#(32) runtime_nhop_ipv4_32;
  } SetNhopReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(2) stats_metadata$flow_map_index;
  } UpdateFlowDupackReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) stats_metadata$flow_map_index;
    Bit#(48) intrinsic_metadata$ingress_global_timestamp;
    Bit#(32) stats_metadata$dummy;
    Bit#(16) tcp$window;
    Bit#(32) tcp$ackNo;
  } UpdateFlowRcvdReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(2) stats_metadata$flow_map_index;
  } UpdateFlowRetx3DupackReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(2) stats_metadata$flow_map_index;
  } UpdateFlowRetxTimeoutReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) stats_metadata$flow_map_index;
    Bit#(48) intrinsic_metadata$ingress_global_timestamp;
    Bit#(32) stats_metadata$dummy;
    Bit#(32) tcp$seqNo;
    Bit#(32) stats_metadata$dummy2;
  } UpdateFlowSentReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(2) stats_metadata$flow_map_index;
    Bit#(48) intrinsic_metadata$ingress_global_timestamp;
  } UseSampleRttReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(2) stats_metadata$flow_map_index;
    Bit#(32) stats_metadata$dummy2;
    Bit#(48) intrinsic_metadata$ingress_global_timestamp;
  } UseSampleRttFirstReqT;
} BBRequest deriving (Bits, Eq, FShow);
typedef union tagged {
  struct {
    PacketInstance pkt;
  } DropRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$sample_rtt_seq;
    Bit#(32) stats_metadata$seqNo;
    Bit#(32) stats_metadata$dupack;
    Bit#(32) stats_metadata$rtt_samples;
    Bit#(32) stats_metadata$ackNo;
    Bit#(32) stats_metadata$senderIP;
    Bit#(32) stats_metadata$mincwnd;
  } GetSenderIpRspT;
  struct {
    PacketInstance pkt;
  } IncreaseMincwndRspT;
  struct {
    PacketInstance pkt;
  } LookupFlowMapRspT;
  struct {
    PacketInstance pkt;
  } LookupFlowMapReverseRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$senderIP;
  } RecordIpRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
  } RewriteMacRspT;
  struct {
    PacketInstance pkt;
  } SampleNewRttRspT;
  struct {
    PacketInstance pkt;
  } SaveSourceIpRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$dstAddr;
  } SetDmacRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ipv4$ttl;
    Bit#(9) standard_metadata$egress_spec;
    Bit#(32) routing_metadata$nhop_ipv4;
  } SetNhopRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
  } UpdateFlowDupackRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
  } UpdateFlowRcvdRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
  } UpdateFlowRetx3DupackRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
  } UpdateFlowRetxTimeoutRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(32) stats_metadata$dummy2;
  } UpdateFlowSentRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(32) stats_metadata$dummy2;
  } UseSampleRttRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) stats_metadata$dummy;
    Bit#(32) stats_metadata$dummy2;
  } UseSampleRttFirstRspT;
} BBResponse deriving (Bits, Eq, FShow);
