import Ethernet::*;
import StructDefines::*;
import Ethernet::*;
import StructDefines::*;
