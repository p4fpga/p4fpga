method Action forward_add_entry(ForwardReqT key, ForwardRspT val);
method Action ipv4_lpm_add_entry(Ipv4LpmReqT key, Ipv4LpmRspT val);
method Action send_frame_add_entry(SendFrameReqT key, SendFrameRspT val);
