method Action forward_table_add_entry(ForwardTableReqT key, ForwardTableRspT val);
method Action table_1_add_entry(Table1ReqT key, Table1RspT val);
method Action table_2_add_entry(Table2ReqT key, Table2RspT val);
method Action table_3_add_entry(Table3ReqT key, Table3RspT val);
method Action table_4_add_entry(Table4ReqT key, Table4RspT val);
method Action table_5_add_entry(Table5ReqT key, Table5RspT val);
method Action table_6_add_entry(Table6ReqT key, Table6RspT val);
method Action table_7_add_entry(Table7ReqT key, Table7RspT val);
