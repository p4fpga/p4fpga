import DefaultValue::*;
import Ethernet::*;
`include "UnionGenerated.bsv"
