method Action forward_add_entry(ForwardReqT key, ForwardRspT val);
method Action ipv4_lpm_add_entry(Ipv4LpmReqT key, Ipv4LpmRspT val);
method Action t_opti_update_add_entry(TOptiUpdateReqT key, TOptiUpdateRspT val);
method Action t_reply_client_add_entry(TReplyClientReqT key, TReplyClientRspT val);
method Action t_req_fix_add_entry(TReqFixReqT key, TReqFixRspT val);
method Action t_req_pass1_add_entry(TReqPass1ReqT key, TReqPass1RspT val);
method Action t_store_update_add_entry(TStoreUpdateReqT key, TStoreUpdateRspT val);
method Action send_frame_add_entry(SendFrameReqT key, SendFrameRspT val);
