method forward_table_add_entry=ingress.forward_table_add_entry;
method test_tbl_add_entry=ingress.test_tbl_add_entry;
