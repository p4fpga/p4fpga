
import BUtils::*;
import BuildVector::*;
import CBus::*;
import ClientServer::*;
import ConfigReg::*;
import Connectable::*;
import DbgDefs::*;
import DefaultValue::*;
import Ethernet::*;
import FIFO::*;
import FIFOF::*;
import FShow::*;
import GetPut::*;
import List::*;
import MIMO::*;
import MatchTable::*;
import PacketBuffer::*;
import Pipe::*;
import PrintTrace::*;
import Register::*;
import SpecialFIFOs::*;
import StmtFSM::*;
import StructGenerated::*;
import TxRx::*;
import Utils::*;
import Vector::*;
typedef union tagged {
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_acl_copy_reason;
    Bit#(1) runtime_acl_copy;
    Bit#(16) runtime_acl_meter_index;
    Bit#(14) runtime_acl_stats_index;
  } AclDenyReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) intrinsic_metadata$ingress_global_tstamp;
    Bit#(32) runtime_session_id;
    Bit#(16) runtime_acl_meter_index;
    Bit#(14) runtime_acl_stats_index;
  } AclMirrorReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_acl_copy_reason;
    Bit#(1) runtime_acl_copy;
    Bit#(16) runtime_acl_meter_index;
    Bit#(14) runtime_acl_stats_index;
  } AclPermitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_acl_copy_reason;
    Bit#(16) runtime_acl_meter_index;
    Bit#(1) runtime_acl_copy;
    Bit#(16) runtime_ecmp_index;
    Bit#(14) runtime_acl_stats_index;
  } AclRedirectEcmpReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_acl_copy_reason;
    Bit#(16) runtime_acl_meter_index;
    Bit#(1) runtime_acl_copy;
    Bit#(16) runtime_nexthop_index;
    Bit#(14) runtime_acl_stats_index;
  } AclRedirectNexthopReqT;
  struct {
    PacketInstance pkt;
  } AclStatsUpdateReqT;
  struct {
    PacketInstance pkt;
    Bit#(3) runtime_cos;
  } ApplyCosMarkingReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_dscp;
  } ApplyDscpMarkingReqT;
  struct {
    PacketInstance pkt;
    Bit#(3) runtime_tc;
  } ApplyTcMarkingReqT;
  struct {
    PacketInstance pkt;
  } ComputeLkpIpv4HashReqT;
  struct {
    PacketInstance pkt;
  } ComputeLkpIpv6HashReqT;
  struct {
    PacketInstance pkt;
  } ComputeLkpNonIpHashReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) hash_metadata$hash2;
  } ComputedOneHashReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) hash_metadata$hash1;
    Bit#(16) hash_metadata$hash2;
  } ComputedTwoHashesReqT;
  struct {
    PacketInstance pkt;
  } CopyToCpuReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_reason_code;
  } CopyToCpuWithReasonReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ingress_metadata$bd;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(9) ingress_metadata$ingress_port;
    Bit#(16) ingress_metadata$ifindex;
    Bit#(16) ethernet$etherType;
  } CpuRxRewriteReqT;
  struct {
    PacketInstance pkt;
  } DecapGenvInnerIpv4ReqT;
  struct {
    PacketInstance pkt;
  } DecapGenvInnerIpv6ReqT;
  struct {
    PacketInstance pkt;
  } DecapGenvInnerNonIpReqT;
  struct {
    PacketInstance pkt;
  } DecapGreInnerIpv4ReqT;
  struct {
    PacketInstance pkt;
  } DecapGreInnerIpv6ReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) gre$proto;
  } DecapGreInnerNonIpReqT;
  struct {
    PacketInstance pkt;
  } DecapInnerIcmpReqT;
  struct {
    PacketInstance pkt;
  } DecapInnerTcpReqT;
  struct {
    PacketInstance pkt;
  } DecapInnerUdpReqT;
  struct {
    PacketInstance pkt;
  } DecapInnerUnknownReqT;
  struct {
    PacketInstance pkt;
  } DecapIpInnerIpv4ReqT;
  struct {
    PacketInstance pkt;
  } DecapIpInnerIpv6ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv4Pop1ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv4Pop2ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv4Pop3ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv6Pop1ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv6Pop2ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv6Pop3ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetNonIpPop1ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetNonIpPop2ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetNonIpPop3ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerIpv4Pop1ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerIpv4Pop2ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerIpv4Pop3ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerIpv6Pop1ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerIpv6Pop2ReqT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerIpv6Pop3ReqT;
  struct {
    PacketInstance pkt;
  } DecapNvgreInnerIpv4ReqT;
  struct {
    PacketInstance pkt;
  } DecapNvgreInnerIpv6ReqT;
  struct {
    PacketInstance pkt;
  } DecapNvgreInnerNonIpReqT;
  struct {
    PacketInstance pkt;
  } DecapVxlanInnerIpv4ReqT;
  struct {
    PacketInstance pkt;
  } DecapVxlanInnerIpv6ReqT;
  struct {
    PacketInstance pkt;
  } DecapVxlanInnerNonIpReqT;
  struct {
    PacketInstance pkt;
  } DmacDropReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_ifindex;
  } DmacHitReqT;
  struct {
    PacketInstance pkt;
  } DmacMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
  } DmacMulticastHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_ecmp_index;
  } DmacRedirectEcmpReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_nexthop_index;
  } DmacRedirectNexthopReqT;
  struct {
    PacketInstance pkt;
  } DropPacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_drop_reason;
  } DropPacketWithReasonReqT;
  struct {
    PacketInstance pkt;
  } DropStatsUpdateReqT;
  struct {
    PacketInstance pkt;
  } EgressFilterCheckReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_session_id;
  } EgressMirrorReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_session_id;
  } EgressMirrorDropReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_ifindex;
  } EgressPortTypeCpuReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_ifindex;
  } EgressPortTypeFabricReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_ifindex;
  } EgressPortTypeNormalReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_reason_code;
  } EgressRedirectToCpuReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) multicast_metadata$mcast_grp;
    Bit#(16) ingress_metadata$bd;
    Bit#(5) tunnel_metadata$ingress_tunnel_type;
    Bit#(1) l3_metadata$routed;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) ingress_metadata$ifindex;
    Bit#(16) ethernet$etherType;
    Bit#(1) l3_metadata$outer_routed;
    Bit#(16) runtime_fabric_mgid;
  } FabricMulticastRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(14) runtime_tunnel_index;
  } FabricRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(5) tunnel_metadata$ingress_tunnel_type;
    Bit#(1) l3_metadata$routed;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) fabric_metadata$dst_port;
    Bit#(16) ethernet$etherType;
    Bit#(1) l3_metadata$outer_routed;
  } FabricUnicastRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_ecmp_index;
  } FibHitEcmpReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_nexthop_index;
  } FibHitNexthopReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(16) runtime_nexthop_index;
  } ForwardMplsReqT;
  struct {
    PacketInstance pkt;
  } GenerateLearnNotifyReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ipv4$totalLen;
  } InnerIpv4IcmpRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ipv4$totalLen;
  } InnerIpv4TcpRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ipv4$totalLen;
  } InnerIpv4UdpRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ipv4$totalLen;
  } InnerIpv4UnknownRewriteReqT;
  struct {
    PacketInstance pkt;
  } InnerIpv6IcmpRewriteReqT;
  struct {
    PacketInstance pkt;
  } InnerIpv6TcpRewriteReqT;
  struct {
    PacketInstance pkt;
  } InnerIpv6UdpRewriteReqT;
  struct {
    PacketInstance pkt;
  } InnerIpv6UnknownRewriteReqT;
  struct {
    PacketInstance pkt;
  } InnerNonIpRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$routed;
    Bit#(14) runtime_tunnel_index;
    Bit#(5) runtime_tunnel_type;
    Bit#(16) runtime_bd;
    Bit#(4) runtime_header_count;
  } InnerReplicaFromRidReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) int_metadata$gpe_int_hdr_len8;
    Bit#(16) int_metadata$insert_byte_cnt;
  } IntAddUpdateVxlanGpeIpv4ReqT;
  struct {
    PacketInstance pkt;
  } IntNoSinkReqT;
  struct {
    PacketInstance pkt;
  } IntResetReqT;
  struct {
    PacketInstance pkt;
  } IntSetEBitReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader0003I0ReqT;
  struct {
    PacketInstance pkt;
    Bit#(19) intrinsic_metadata$enq_qdepth;
  } IntSetHeader0003I1ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) intrinsic_metadata$deq_timedelta;
    Bit#(32) int_metadata$switch_id;
  } IntSetHeader0003I10ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) intrinsic_metadata$deq_timedelta;
    Bit#(19) intrinsic_metadata$enq_qdepth;
    Bit#(32) int_metadata$switch_id;
  } IntSetHeader0003I11ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) int_metadata$switch_id;
    Bit#(16) ingress_metadata$ifindex;
  } IntSetHeader0003I12ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) int_metadata$switch_id;
    Bit#(19) intrinsic_metadata$enq_qdepth;
    Bit#(16) ingress_metadata$ifindex;
  } IntSetHeader0003I13ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) intrinsic_metadata$deq_timedelta;
    Bit#(16) ingress_metadata$ifindex;
    Bit#(32) int_metadata$switch_id;
  } IntSetHeader0003I14ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) intrinsic_metadata$deq_timedelta;
    Bit#(19) intrinsic_metadata$enq_qdepth;
    Bit#(16) ingress_metadata$ifindex;
    Bit#(32) int_metadata$switch_id;
  } IntSetHeader0003I15ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) intrinsic_metadata$deq_timedelta;
  } IntSetHeader0003I2ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) intrinsic_metadata$deq_timedelta;
    Bit#(19) intrinsic_metadata$enq_qdepth;
  } IntSetHeader0003I3ReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ingress_metadata$ifindex;
  } IntSetHeader0003I4ReqT;
  struct {
    PacketInstance pkt;
    Bit#(19) intrinsic_metadata$enq_qdepth;
    Bit#(16) ingress_metadata$ifindex;
  } IntSetHeader0003I5ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) intrinsic_metadata$deq_timedelta;
    Bit#(16) ingress_metadata$ifindex;
  } IntSetHeader0003I6ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) intrinsic_metadata$deq_timedelta;
    Bit#(19) intrinsic_metadata$enq_qdepth;
    Bit#(16) ingress_metadata$ifindex;
  } IntSetHeader0003I7ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) int_metadata$switch_id;
  } IntSetHeader0003I8ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) int_metadata$switch_id;
    Bit#(19) intrinsic_metadata$enq_qdepth;
  } IntSetHeader0003I9ReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader0407I0ReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader0407I1ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
  } IntSetHeader0407I10ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
  } IntSetHeader0407I11ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
    Bit#(9) standard_metadata$egress_port;
  } IntSetHeader0407I12ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
    Bit#(9) standard_metadata$egress_port;
  } IntSetHeader0407I13ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
    Bit#(9) standard_metadata$egress_port;
  } IntSetHeader0407I14ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
    Bit#(9) standard_metadata$egress_port;
  } IntSetHeader0407I15ReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader0407I2ReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader0407I3ReqT;
  struct {
    PacketInstance pkt;
    Bit#(9) standard_metadata$egress_port;
  } IntSetHeader0407I4ReqT;
  struct {
    PacketInstance pkt;
    Bit#(9) standard_metadata$egress_port;
  } IntSetHeader0407I5ReqT;
  struct {
    PacketInstance pkt;
    Bit#(9) standard_metadata$egress_port;
  } IntSetHeader0407I6ReqT;
  struct {
    PacketInstance pkt;
    Bit#(9) standard_metadata$egress_port;
  } IntSetHeader0407I7ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
  } IntSetHeader0407I8ReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
  } IntSetHeader0407I9ReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader0BosReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader1BosReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader2BosReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader3BosReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader4BosReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader5BosReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader6BosReqT;
  struct {
    PacketInstance pkt;
  } IntSetHeader7BosReqT;
  struct {
    PacketInstance pkt;
  } IntSetNoSrcReqT;
  struct {
    PacketInstance pkt;
  } IntSetSrcReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_mirror_id;
  } IntSinkGpeReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) vxlan_gpe_int_header$next_proto;
  } IntSinkUpdateVxlanGpeV4ReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_total_words;
    Bit#(32) runtime_switch_id;
    Bit#(4) runtime_ins_mask0003;
    Bit#(16) runtime_ins_byte_cnt;
    Bit#(5) runtime_ins_cnt;
    Bit#(8) runtime_hop_cnt;
    Bit#(4) runtime_ins_mask0407;
  } IntSrcReqT;
  struct {
    PacketInstance pkt;
    Bit#(5) int_header$ins_cnt;
    Bit#(32) runtime_switch_id;
  } IntTransitReqT;
  struct {
    PacketInstance pkt;
  } IntUpdateTotalHopCntReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) int_metadata$gpe_int_hdr_len8;
    Bit#(16) int_metadata$insert_byte_cnt;
  } IntUpdateVxlanGpeIpv4ReqT;
  struct {
    PacketInstance pkt;
  } IpsgMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
    Bit#(16) i2e_metadata$mirror_session_id;
  } Ipv4ErspanT3RewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) hash_metadata$entropy_hash;
    Bit#(24) tunnel_metadata$vnid;
  } Ipv4GenvRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } Ipv4GreRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
  } Ipv4IpRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_l3_mtu;
  } Ipv4MtuCheckReqT;
  struct {
    PacketInstance pkt;
  } Ipv4MulticastRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(24) tunnel_metadata$vnid;
  } Ipv4NvgreRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(32) ipv4$srcAddr;
    Bit#(32) ipv4$dstAddr;
    Bit#(16) l3_metadata$lkp_outer_l4_dport;
    Bit#(8) ipv4$protocol;
    Bit#(16) l3_metadata$lkp_outer_l4_sport;
  } Ipv4OverFabricReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$lkp_outer_l4_dport;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(32) ipv4$srcAddr;
    Bit#(32) ipv4$dstAddr;
    Bit#(8) ipv4$ttl;
    Bit#(8) ipv4$protocol;
    Bit#(16) l3_metadata$lkp_outer_l4_sport;
  } Ipv4TunnelLookupMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) egress_metadata$mac_da;
  } Ipv4UnicastRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) ipv4_metadata$ipv4_urpf_mode;
    Bit#(16) runtime_urpf_bd_group;
  } Ipv4UrpfHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) hash_metadata$entropy_hash;
    Bit#(24) tunnel_metadata$vnid;
  } Ipv4VxlanRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
    Bit#(16) i2e_metadata$mirror_session_id;
  } Ipv6ErspanT3RewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) hash_metadata$entropy_hash;
    Bit#(24) tunnel_metadata$vnid;
  } Ipv6GenvRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } Ipv6GreRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
    Bit#(16) egress_metadata$payload_length;
  } Ipv6IpRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_l3_mtu;
  } Ipv6MtuCheckReqT;
  struct {
    PacketInstance pkt;
  } Ipv6MulticastRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(24) tunnel_metadata$vnid;
  } Ipv6NvgreRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(128) ipv6$srcAddr;
    Bit#(16) l3_metadata$lkp_outer_l4_dport;
    Bit#(128) ipv6$dstAddr;
    Bit#(8) ipv6$nextHdr;
    Bit#(16) l3_metadata$lkp_outer_l4_sport;
  } Ipv6OverFabricReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(128) ipv6$srcAddr;
    Bit#(16) l3_metadata$lkp_outer_l4_dport;
    Bit#(128) ipv6$dstAddr;
    Bit#(8) ipv6$hopLimit;
    Bit#(8) ipv6$nextHdr;
    Bit#(16) l3_metadata$lkp_outer_l4_sport;
  } Ipv6TunnelLookupMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) egress_metadata$mac_da;
  } Ipv6UnicastRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) ipv6_metadata$ipv6_urpf_mode;
    Bit#(16) runtime_urpf_bd_group;
  } Ipv6UrpfHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) hash_metadata$entropy_hash;
    Bit#(24) tunnel_metadata$vnid;
  } Ipv6VxlanRewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_drop_reason;
  } MalformedOuterEthernetPacketReqT;
  struct {
    PacketInstance pkt;
  } MeterDenyReqT;
  struct {
    PacketInstance pkt;
  } MeterPermitReqT;
  struct {
    PacketInstance pkt;
  } MplsEthernetPush1RewriteReqT;
  struct {
    PacketInstance pkt;
  } MplsEthernetPush2RewriteReqT;
  struct {
    PacketInstance pkt;
  } MplsEthernetPush3RewriteReqT;
  struct {
    PacketInstance pkt;
  } MplsIpPush1RewriteReqT;
  struct {
    PacketInstance pkt;
  } MplsIpPush2RewriteReqT;
  struct {
    PacketInstance pkt;
  } MplsIpPush3RewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) egress_metadata$mac_da;
  } MplsRewriteReqT;
  struct {
    PacketInstance pkt;
  } MtuMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
  } MulticastBridgeSGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
  } MulticastBridgeStarGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
    Bit#(16) runtime_mcast_rpf_group;
  } MulticastRouteBidirStarGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
    Bit#(16) runtime_mcast_rpf_group;
  } MulticastRouteSGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
    Bit#(16) runtime_mcast_rpf_group;
  } MulticastRouteSmStarGHitReqT;
  struct {
    PacketInstance pkt;
  } MulticastRouteStarGMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_session_id;
  } NegativeMirrorReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(16) ethernet$etherType;
  } NonIpOverFabricReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
  } NonIpTunnelLookupMissReqT;
  struct {
    PacketInstance pkt;
  } NopReqT;
  struct {
    PacketInstance pkt;
  } OnMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
  } OuterMulticastBridgeSGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
  } OuterMulticastBridgeStarGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
    Bit#(16) runtime_mcast_rpf_group;
  } OuterMulticastRouteBidirStarGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
    Bit#(16) runtime_mcast_rpf_group;
  } OuterMulticastRouteSGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
    Bit#(16) runtime_mcast_rpf_group;
  } OuterMulticastRouteSmStarGHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$outer_routed;
    Bit#(14) runtime_tunnel_index;
    Bit#(5) runtime_tunnel_type;
    Bit#(16) runtime_bd;
    Bit#(4) runtime_header_count;
  } OuterReplicaFromRidReqT;
  struct {
    PacketInstance pkt;
  } OuterRmacHitReqT;
  struct {
    PacketInstance pkt;
  } PortVlanMappingMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) runtime_acl_copy;
    Bit#(16) runtime_acl_copy_reason;
    Bit#(14) runtime_acl_stats_index;
  } RaclDenyReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) runtime_acl_copy;
    Bit#(16) runtime_acl_copy_reason;
    Bit#(14) runtime_acl_stats_index;
  } RaclPermitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_acl_copy_reason;
    Bit#(1) runtime_acl_copy;
    Bit#(16) runtime_ecmp_index;
    Bit#(14) runtime_acl_stats_index;
  } RaclRedirectEcmpReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_acl_copy_reason;
    Bit#(1) runtime_acl_copy;
    Bit#(16) runtime_nexthop_index;
    Bit#(14) runtime_acl_stats_index;
  } RaclRedirectNexthopReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_reason_code;
  } RedirectToCpuReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) vlan_tag_1$etherType;
  } RemoveVlanDoubleTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) vlan_tag_0$etherType;
  } RemoveVlanSingleTaggedReqT;
  struct {
    PacketInstance pkt;
  } RewriteIpv4MulticastReqT;
  struct {
    PacketInstance pkt;
  } RewriteIpv6MulticastReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) runtime_smac;
  } RewriteSmacReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) runtime_dmac;
  } RewriteTunnelDmacReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_ip;
  } RewriteTunnelIpv4DstReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_ip;
  } RewriteTunnelIpv4SrcReqT;
  struct {
    PacketInstance pkt;
    Bit#(128) runtime_ip;
  } RewriteTunnelIpv6DstReqT;
  struct {
    PacketInstance pkt;
    Bit#(128) runtime_ip;
  } RewriteTunnelIpv6SrcReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) runtime_smac;
  } RewriteTunnelSmacReqT;
  struct {
    PacketInstance pkt;
  } RmacHitReqT;
  struct {
    PacketInstance pkt;
  } RmacMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) acl_metadata$acl_nexthop;
    Bit#(1) acl_metadata$acl_nexthop_type;
  } SetAclRedirectActionReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_mc_index;
  } SetBdFloodMcIndexReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) runtime_ipv4_multicast_enabled;
    Bit#(1) runtime_igmp_snooping_enabled;
    Bit#(16) runtime_ipv6_mcast_key;
    Bit#(16) runtime_mrpf_group;
    Bit#(1) runtime_ipv4_mcast_key_type;
    Bit#(1) runtime_mld_snooping_enabled;
    Bit#(1) runtime_ipv6_multicast_enabled;
    Bit#(16) runtime_stats_idx;
    Bit#(2) runtime_ipv6_urpf_mode;
    Bit#(2) runtime_ipv4_urpf_mode;
    Bit#(16) runtime_ipv4_mcast_key;
    Bit#(16) runtime_bd;
    Bit#(16) runtime_vrf;
    Bit#(1) runtime_learning_enabled;
    Bit#(1) runtime_ipv6_unicast_enabled;
    Bit#(16) runtime_bd_label;
    Bit#(1) runtime_ipv6_mcast_key_type;
    Bit#(10) runtime_rmac_group;
    Bit#(1) runtime_ipv4_unicast_enabled;
    Bit#(10) runtime_stp_group;
  } SetBdPropertiesReqT;
  struct {
    PacketInstance pkt;
  } SetBroadcastReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ingress_metadata$ifindex;
    Bit#(48) intrinsic_metadata$ingress_global_tstamp;
    Bit#(9) standard_metadata$ingress_port;
    Bit#(1) runtime_enable_dod;
  } SetConfigParametersReqT;
  struct {
    PacketInstance pkt;
  } SetCpuRedirectActionReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_bd;
    Bit#(16) runtime_nhop_index;
    Bit#(16) runtime_ifindex;
    Bit#(1) runtime_tunnel;
  } SetEcmpNexthopDetailsReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_uuc_mc_index;
    Bit#(16) runtime_nhop_index;
    Bit#(16) runtime_bd;
  } SetEcmpNexthopDetailsForPostRoutedFloodReqT;
  struct {
    PacketInstance pkt;
    Bit#(9) runtime_smac_idx;
  } SetEgressBdPropertiesReqT;
  struct {
    PacketInstance pkt;
  } SetEgressFilterDropReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
    Bit#(12) runtime_c_tag;
    Bit#(12) runtime_s_tag;
  } SetEgressPacketVlanDoubleTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
    Bit#(12) runtime_vlan_id;
  } SetEgressPacketVlanTaggedReqT;
  struct {
    PacketInstance pkt;
  } SetEgressPacketVlanUntaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(24) runtime_vnid;
  } SetEgressTunnelVniReqT;
  struct {
    PacketInstance pkt;
    Bit#(9) runtime_port;
  } SetFabricLagPortReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } SetFabricMulticastReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$fib_nexthop;
    Bit#(1) l3_metadata$fib_nexthop_type;
  } SetFibRedirectActionReqT;
  struct {
    PacketInstance pkt;
    Bit#(2) runtime_port_type;
    Bit#(16) runtime_ifindex;
  } SetIfindexReqT;
  struct {
    PacketInstance pkt;
  } SetIngressIfindexPropertiesReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_if_label;
  } SetIngressPortPropertiesReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) l2_metadata$l2_nexthop;
    Bit#(1) l2_metadata$l2_nexthop_type;
  } SetL2RedirectActionReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ingress_metadata$bd;
  } SetL2RewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ingress_metadata$bd;
    Bit#(14) runtime_tunnel_index;
    Bit#(5) runtime_tunnel_type;
  } SetL2RewriteWithTunnelReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) runtime_dmac;
    Bit#(16) runtime_bd;
    Bit#(8) runtime_mtu_index;
  } SetL3RewriteReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) runtime_dmac;
    Bit#(14) runtime_tunnel_index;
    Bit#(16) runtime_bd;
    Bit#(5) runtime_tunnel_type;
  } SetL3RewriteWithTunnelReqT;
  struct {
    PacketInstance pkt;
  } SetLagMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(9) runtime_port;
  } SetLagPortReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_device;
    Bit#(16) runtime_port;
  } SetLagRemotePortReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_drop_reason;
  } SetMalformedOuterIpv4PacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_drop_reason;
  } SetMalformedOuterIpv6PacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_drop_reason;
  } SetMalformedPacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_bd;
  } SetMirrorBdReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_nhop_idx;
  } SetMirrorNhopReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$routed;
    Bit#(16) ingress_metadata$bd;
    Bit#(14) runtime_tunnel_index;
    Bit#(4) runtime_header_count;
  } SetMplsPushRewriteL2ReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$routed;
    Bit#(48) runtime_dmac;
    Bit#(14) runtime_tunnel_index;
    Bit#(16) runtime_bd;
    Bit#(4) runtime_header_count;
  } SetMplsPushRewriteL3ReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_ttl1;
    Bit#(3) runtime_exp1;
    Bit#(20) runtime_label1;
    Bit#(14) runtime_dmac_idx;
    Bit#(9) runtime_smac_idx;
  } SetMplsRewritePush1ReqT;
  struct {
    PacketInstance pkt;
    Bit#(3) runtime_exp1;
    Bit#(8) runtime_ttl2;
    Bit#(9) runtime_smac_idx;
    Bit#(8) runtime_ttl1;
    Bit#(20) runtime_label2;
    Bit#(3) runtime_exp2;
    Bit#(20) runtime_label1;
    Bit#(14) runtime_dmac_idx;
  } SetMplsRewritePush2ReqT;
  struct {
    PacketInstance pkt;
    Bit#(3) runtime_exp3;
    Bit#(3) runtime_exp1;
    Bit#(8) runtime_ttl2;
    Bit#(20) runtime_label3;
    Bit#(8) runtime_ttl1;
    Bit#(20) runtime_label2;
    Bit#(3) runtime_exp2;
    Bit#(20) runtime_label1;
    Bit#(9) runtime_smac_idx;
    Bit#(8) runtime_ttl3;
    Bit#(14) runtime_dmac_idx;
  } SetMplsRewritePush3ReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$routed;
    Bit#(16) ingress_metadata$bd;
    Bit#(14) runtime_tunnel_index;
    Bit#(20) runtime_label;
    Bit#(4) runtime_header_count;
  } SetMplsSwapPushRewriteL2ReqT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$routed;
    Bit#(48) runtime_dmac;
    Bit#(14) runtime_tunnel_index;
    Bit#(20) runtime_label;
    Bit#(16) runtime_bd;
    Bit#(4) runtime_header_count;
  } SetMplsSwapPushRewriteL3ReqT;
  struct {
    PacketInstance pkt;
  } SetMulticastReqT;
  struct {
    PacketInstance pkt;
  } SetMulticastAndIpv6SrcIsLinkLocalReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) multicast_metadata$multicast_bridge_mc_index;
  } SetMulticastBridgeActionReqT;
  struct {
    PacketInstance pkt;
  } SetMulticastDropReqT;
  struct {
    PacketInstance pkt;
  } SetMulticastFloodReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) multicast_metadata$multicast_route_mc_index;
  } SetMulticastRouteActionReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_bd;
    Bit#(1) runtime_tunnel;
    Bit#(16) runtime_ifindex;
  } SetNexthopDetailsReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_uuc_mc_index;
    Bit#(16) runtime_bd;
  } SetNexthopDetailsForPostRoutedFloodReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) acl_metadata$racl_nexthop;
    Bit#(1) acl_metadata$racl_nexthop_type;
  } SetRaclRedirectActionReqT;
  struct {
    PacketInstance pkt;
  } SetReplicaCopyBridgedReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_meter_idx;
  } SetStormControlMeterReqT;
  struct {
    PacketInstance pkt;
    Bit#(3) runtime_stp_state;
  } SetStpStateReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_outer_bd;
    Bit#(9) runtime_sip_index;
    Bit#(14) runtime_dip_index;
    Bit#(14) runtime_dmac_idx;
    Bit#(9) runtime_smac_idx;
  } SetTunnelRewriteDetailsReqT;
  struct {
    PacketInstance pkt;
  } SetTunnelTerminationFlagReqT;
  struct {
    PacketInstance pkt;
    Bit#(24) runtime_tunnel_vni;
  } SetTunnelVniAndTerminationFlagReqT;
  struct {
    PacketInstance pkt;
  } SetUnicastReqT;
  struct {
    PacketInstance pkt;
  } SetUnicastAndIpv6SrcIsLinkLocalReqT;
  struct {
    PacketInstance pkt;
    Bit#(3) mpls0$exp;
    Bit#(20) mpls0$label;
  } SetValidMplsLabel1ReqT;
  struct {
    PacketInstance pkt;
    Bit#(20) mpls1$label;
    Bit#(3) mpls1$exp;
  } SetValidMplsLabel2ReqT;
  struct {
    PacketInstance pkt;
    Bit#(20) mpls2$label;
    Bit#(3) mpls2$exp;
  } SetValidMplsLabel3ReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) vlan_tag_1$etherType;
  } SetValidOuterBroadcastPacketDoubleTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } SetValidOuterBroadcastPacketQinqTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) vlan_tag_0$etherType;
  } SetValidOuterBroadcastPacketSingleTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } SetValidOuterBroadcastPacketUntaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) ipv4$diffserv;
    Bit#(4) ipv4$version;
  } SetValidOuterIpv4PacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(4) ipv6$version;
    Bit#(8) ipv6$trafficClass;
  } SetValidOuterIpv6PacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) vlan_tag_1$etherType;
  } SetValidOuterMulticastPacketDoubleTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } SetValidOuterMulticastPacketQinqTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) vlan_tag_0$etherType;
  } SetValidOuterMulticastPacketSingleTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } SetValidOuterMulticastPacketUntaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) vlan_tag_1$etherType;
  } SetValidOuterUnicastPacketDoubleTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } SetValidOuterUnicastPacketQinqTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) vlan_tag_0$etherType;
  } SetValidOuterUnicastPacketSingleTaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } SetValidOuterUnicastPacketUntaggedReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_sflow_i2e_mirror_id;
    Bit#(16) runtime_reason_code;
  } SflowIngPktToCpuReqT;
  struct {
    PacketInstance pkt;
    Bit#(32) runtime_rate_thr;
    Bit#(16) runtime_session_id;
  } SflowIngSessionEnableReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) sflow_metadata$sflow_session_id;
  } SflowPktToCpuReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_ifindex;
  } SmacHitReqT;
  struct {
    PacketInstance pkt;
  } SmacMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_ifindex;
  } SrcVtepHitReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) fabric_header$dstPortOrGroup;
  } SwitchFabricMulticastPacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_header$dstDevice;
    Bit#(16) fabric_header$dstPortOrGroup;
  } SwitchFabricUnicastPacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) fabric_payload_header$etherType;
    Bit#(1) fabric_header_cpu$txBypass;
    Bit#(16) fabric_header$dstPortOrGroup;
  } TerminateCpuPacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) inner_ethernet$etherType;
    Bit#(5) runtime_tunnel_type;
    Bit#(16) runtime_bd;
  } TerminateEomplsReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) fabric_payload_header$etherType;
    Bit#(1) fabric_header_multicast$tunnelTerminate;
    Bit#(1) fabric_header_multicast$outerRouted;
    Bit#(5) fabric_header_multicast$ingressTunnelType;
    Bit#(16) fabric_header_multicast$mcastGrp;
    Bit#(1) fabric_header_multicast$routed;
  } TerminateFabricMulticastPacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) fabric_header_unicast$nexthopIndex;
    Bit#(1) fabric_header_unicast$routed;
    Bit#(1) fabric_header_unicast$tunnelTerminate;
    Bit#(16) fabric_payload_header$etherType;
    Bit#(1) fabric_header_unicast$outerRouted;
    Bit#(5) fabric_header_unicast$ingressTunnelType;
    Bit#(16) fabric_header$dstPortOrGroup;
  } TerminateFabricUnicastPacketReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) inner_ipv4$diffserv;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(16) inner_ethernet$etherType;
    Bit#(4) inner_ipv4$version;
    Bit#(5) runtime_tunnel_type;
    Bit#(16) runtime_vrf;
  } TerminateIpv4OverMplsReqT;
  struct {
    PacketInstance pkt;
    Bit#(4) inner_ipv6$version;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(16) inner_ethernet$etherType;
    Bit#(8) inner_ipv6$trafficClass;
    Bit#(5) runtime_tunnel_type;
    Bit#(16) runtime_vrf;
  } TerminateIpv6OverMplsReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(16) runtime_ifindex;
  } TerminatePwReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(4) inner_ipv4$version;
    Bit#(16) inner_ethernet$etherType;
    Bit#(8) inner_ipv4$diffserv;
    Bit#(1) runtime_ipv4_multicast_enabled;
    Bit#(1) runtime_igmp_snooping_enabled;
    Bit#(16) runtime_mrpf_group;
    Bit#(16) runtime_stats_idx;
    Bit#(2) runtime_ipv4_urpf_mode;
    Bit#(16) runtime_bd;
    Bit#(16) runtime_vrf;
    Bit#(16) runtime_bd_label;
    Bit#(10) runtime_rmac_group;
    Bit#(1) runtime_ipv4_unicast_enabled;
  } TerminateTunnelInnerEthernetIpv4ReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(8) inner_ipv6$trafficClass;
    Bit#(16) inner_ethernet$etherType;
    Bit#(4) inner_ipv6$version;
    Bit#(16) runtime_mrpf_group;
    Bit#(1) runtime_mld_snooping_enabled;
    Bit#(1) runtime_ipv6_multicast_enabled;
    Bit#(16) runtime_stats_idx;
    Bit#(2) runtime_ipv6_urpf_mode;
    Bit#(16) runtime_bd;
    Bit#(16) runtime_vrf;
    Bit#(1) runtime_ipv6_unicast_enabled;
    Bit#(16) runtime_bd_label;
    Bit#(10) runtime_rmac_group;
  } TerminateTunnelInnerEthernetIpv6ReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(8) inner_ipv4$diffserv;
    Bit#(4) inner_ipv4$version;
    Bit#(1) runtime_ipv4_multicast_enabled;
    Bit#(16) runtime_mrpf_group;
    Bit#(2) runtime_ipv4_urpf_mode;
    Bit#(16) runtime_vrf;
    Bit#(10) runtime_rmac_group;
    Bit#(1) runtime_ipv4_unicast_enabled;
  } TerminateTunnelInnerIpv4ReqT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
    Bit#(48) ethernet$dstAddr;
    Bit#(128) inner_ipv6$dstAddr;
    Bit#(128) inner_ipv6$srcAddr;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(8) inner_ipv6$trafficClass;
    Bit#(4) inner_ipv6$version;
    Bit#(16) runtime_mrpf_group;
    Bit#(1) runtime_ipv6_multicast_enabled;
    Bit#(2) runtime_ipv6_urpf_mode;
    Bit#(16) runtime_vrf;
    Bit#(1) runtime_ipv6_unicast_enabled;
    Bit#(10) runtime_rmac_group;
  } TerminateTunnelInnerIpv6ReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) inner_ethernet$etherType;
    Bit#(16) runtime_bd_label;
    Bit#(16) runtime_bd;
    Bit#(16) runtime_stats_idx;
  } TerminateTunnelInnerNonIpReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) inner_ethernet$etherType;
    Bit#(5) runtime_tunnel_type;
    Bit#(16) runtime_bd;
  } TerminateVplsReqT;
  struct {
    PacketInstance pkt;
  } TunnelLookupMissReqT;
  struct {
    PacketInstance pkt;
    Bit#(16) runtime_l3_mtu;
  } TunnelMtuCheckReqT;
  struct {
    PacketInstance pkt;
  } TunnelMtuMissReqT;
  struct {
    PacketInstance pkt;
  } UpdateIngressBdStatsReqT;
  struct {
    PacketInstance pkt;
  } UrpfBdMissReqT;
  struct {
    PacketInstance pkt;
  } UrpfMissReqT;
} BBRequest deriving (Bits, Eq, FShow);
typedef union tagged {
  struct {
    PacketInstance pkt;
    Bit#(1) acl_metadata$acl_deny;
    Bit#(14) acl_metadata$acl_stats_index;
    Bit#(16) meter_metadata$meter_index;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(1) acl_metadata$acl_copy;
  } AclDenyRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) i2e_metadata$ingress_tstamp;
    Bit#(14) acl_metadata$acl_stats_index;
    Bit#(16) meter_metadata$meter_index;
    Bit#(16) i2e_metadata$mirror_session_id;
  } AclMirrorRspT;
  struct {
    PacketInstance pkt;
    Bit#(14) acl_metadata$acl_stats_index;
    Bit#(16) meter_metadata$meter_index;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(1) acl_metadata$acl_copy;
  } AclPermitRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) meter_metadata$meter_index;
    Bit#(14) acl_metadata$acl_stats_index;
    Bit#(1) acl_metadata$acl_redirect;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(16) acl_metadata$acl_nexthop;
    Bit#(1) acl_metadata$acl_copy;
    Bit#(1) acl_metadata$acl_nexthop_type;
  } AclRedirectEcmpRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) meter_metadata$meter_index;
    Bit#(14) acl_metadata$acl_stats_index;
    Bit#(1) acl_metadata$acl_redirect;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(16) acl_metadata$acl_nexthop;
    Bit#(1) acl_metadata$acl_copy;
    Bit#(1) acl_metadata$acl_nexthop_type;
  } AclRedirectNexthopRspT;
  struct {
    PacketInstance pkt;
  } AclStatsUpdateRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) qos_metadata$marked_cos;
  } ApplyCosMarkingRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) qos_metadata$marked_dscp;
  } ApplyDscpMarkingRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) qos_metadata$marked_exp;
  } ApplyTcMarkingRspT;
  struct {
    PacketInstance pkt;
  } ComputeLkpIpv4HashRspT;
  struct {
    PacketInstance pkt;
  } ComputeLkpIpv6HashRspT;
  struct {
    PacketInstance pkt;
  } ComputeLkpNonIpHashRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) hash_metadata$entropy_hash;
    Bit#(13) intrinsic_metadata$mcast_hash;
    Bit#(16) hash_metadata$hash1;
  } ComputedOneHashRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) hash_metadata$entropy_hash;
    Bit#(13) intrinsic_metadata$mcast_hash;
  } ComputedTwoHashesRspT;
  struct {
    PacketInstance pkt;
  } CopyToCpuRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) fabric_metadata$reason_code;
  } CopyToCpuWithReasonRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) fabric_header$packetType;
    Bit#(16) fabric_header_cpu$reasonCode;
    Bit#(16) fabric_header_cpu$ingressPort;
    Bit#(16) fabric_header_cpu$ingressIfindex;
    Bit#(16) fabric_payload_header$etherType;
    Bit#(16) fabric_header_cpu$ingressBd;
    Bit#(2) fabric_header$headerVersion;
    Bit#(2) fabric_header$packetVersion;
    Bit#(16) ethernet$etherType;
    Bit#(1) fabric_header$pad1;
  } CpuRxRewriteRspT;
  struct {
    PacketInstance pkt;
  } DecapGenvInnerIpv4RspT;
  struct {
    PacketInstance pkt;
  } DecapGenvInnerIpv6RspT;
  struct {
    PacketInstance pkt;
  } DecapGenvInnerNonIpRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapGreInnerIpv4RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapGreInnerIpv6RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapGreInnerNonIpRspT;
  struct {
    PacketInstance pkt;
  } DecapInnerIcmpRspT;
  struct {
    PacketInstance pkt;
  } DecapInnerTcpRspT;
  struct {
    PacketInstance pkt;
  } DecapInnerUdpRspT;
  struct {
    PacketInstance pkt;
  } DecapInnerUnknownRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapIpInnerIpv4RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapIpInnerIpv6RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv4Pop1RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv4Pop2RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv4Pop3RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv6Pop1RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv6Pop2RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetIpv6Pop3RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetNonIpPop1RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetNonIpPop2RspT;
  struct {
    PacketInstance pkt;
  } DecapMplsInnerEthernetNonIpPop3RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapMplsInnerIpv4Pop1RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapMplsInnerIpv4Pop2RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapMplsInnerIpv4Pop3RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapMplsInnerIpv6Pop1RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapMplsInnerIpv6Pop2RspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } DecapMplsInnerIpv6Pop3RspT;
  struct {
    PacketInstance pkt;
  } DecapNvgreInnerIpv4RspT;
  struct {
    PacketInstance pkt;
  } DecapNvgreInnerIpv6RspT;
  struct {
    PacketInstance pkt;
  } DecapNvgreInnerNonIpRspT;
  struct {
    PacketInstance pkt;
  } DecapVxlanInnerIpv4RspT;
  struct {
    PacketInstance pkt;
  } DecapVxlanInnerIpv6RspT;
  struct {
    PacketInstance pkt;
  } DecapVxlanInnerNonIpRspT;
  struct {
    PacketInstance pkt;
  } DmacDropRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ingress_metadata$egress_ifindex;
  } DmacHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) ingress_metadata$egress_ifindex;
  } DmacMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } DmacMulticastHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l2_metadata$l2_redirect;
    Bit#(16) l2_metadata$l2_nexthop;
    Bit#(1) l2_metadata$l2_nexthop_type;
  } DmacRedirectEcmpRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l2_metadata$l2_redirect;
    Bit#(16) l2_metadata$l2_nexthop;
    Bit#(1) l2_metadata$l2_nexthop_type;
  } DmacRedirectNexthopRspT;
  struct {
    PacketInstance pkt;
  } DropPacketRspT;
  struct {
    PacketInstance pkt;
  } DropPacketWithReasonRspT;
  struct {
    PacketInstance pkt;
  } DropStatsUpdateRspT;
  struct {
    PacketInstance pkt;
  } EgressFilterCheckRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) i2e_metadata$mirror_session_id;
  } EgressMirrorRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) i2e_metadata$mirror_session_id;
  } EgressMirrorDropRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$ifindex;
    Bit#(2) egress_metadata$port_type;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
  } EgressPortTypeCpuRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$ifindex;
    Bit#(2) egress_metadata$port_type;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
  } EgressPortTypeFabricRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$ifindex;
    Bit#(2) egress_metadata$port_type;
  } EgressPortTypeNormalRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) fabric_metadata$reason_code;
  } EgressRedirectToCpuRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) fabric_header$packetType;
    Bit#(1) fabric_header_multicast$tunnelTerminate;
    Bit#(1) fabric_header_multicast$routed;
    Bit#(5) fabric_header_multicast$ingressTunnelType;
    Bit#(8) fabric_header$dstDevice;
    Bit#(1) fabric_header_multicast$outerRouted;
    Bit#(16) fabric_header_multicast$ingressIfindex;
    Bit#(16) fabric_header$dstPortOrGroup;
    Bit#(16) fabric_payload_header$etherType;
    Bit#(16) fabric_header_multicast$ingressBd;
    Bit#(16) fabric_header_multicast$mcastGrp;
    Bit#(1) fabric_header$pad1;
    Bit#(2) fabric_header$packetVersion;
    Bit#(16) ethernet$etherType;
    Bit#(2) fabric_header$headerVersion;
  } FabricMulticastRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(14) tunnel_metadata$tunnel_index;
  } FabricRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) fabric_header$packetType;
    Bit#(1) fabric_header_unicast$outerRouted;
    Bit#(1) fabric_header_unicast$tunnelTerminate;
    Bit#(16) fabric_payload_header$etherType;
    Bit#(8) fabric_header$dstDevice;
    Bit#(5) fabric_header_unicast$ingressTunnelType;
    Bit#(16) fabric_header$dstPortOrGroup;
    Bit#(16) fabric_header_unicast$nexthopIndex;
    Bit#(1) fabric_header_unicast$routed;
    Bit#(1) fabric_header$pad1;
    Bit#(2) fabric_header$packetVersion;
    Bit#(16) ethernet$etherType;
    Bit#(2) fabric_header$headerVersion;
  } FabricUnicastRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$fib_nexthop;
    Bit#(1) l3_metadata$fib_hit;
    Bit#(1) l3_metadata$fib_nexthop_type;
  } FibHitEcmpRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$fib_nexthop;
    Bit#(1) l3_metadata$fib_hit;
    Bit#(1) l3_metadata$fib_nexthop_type;
  } FibHitNexthopRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(16) l3_metadata$fib_nexthop;
    Bit#(1) l3_metadata$fib_hit;
    Bit#(1) l3_metadata$fib_nexthop_type;
    Bit#(48) l2_metadata$lkp_mac_da;
  } ForwardMplsRspT;
  struct {
    PacketInstance pkt;
  } GenerateLearnNotifyRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
    Bit#(16) egress_metadata$payload_length;
  } InnerIpv4IcmpRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
    Bit#(16) egress_metadata$payload_length;
  } InnerIpv4TcpRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
    Bit#(16) egress_metadata$payload_length;
  } InnerIpv4UdpRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
    Bit#(16) egress_metadata$payload_length;
  } InnerIpv4UnknownRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
  } InnerIpv6IcmpRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
  } InnerIpv6TcpRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
  } InnerIpv6UdpRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) tunnel_metadata$inner_ip_proto;
  } InnerIpv6UnknownRewriteRspT;
  struct {
    PacketInstance pkt;
  } InnerNonIpRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) multicast_metadata$replica;
    Bit#(1) multicast_metadata$inner_replica;
    Bit#(4) tunnel_metadata$egress_header_count;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
    Bit#(16) egress_metadata$bd;
    Bit#(14) tunnel_metadata$tunnel_index;
    Bit#(1) egress_metadata$routed;
  } InnerReplicaFromRidRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) vxlan_gpe$next_proto;
    Bit#(8) vxlan_gpe_int_header$len;
    Bit#(8) vxlan_gpe_int_header$next_proto;
    Bit#(8) vxlan_gpe_int_header$int_type;
    Bit#(16) udp$length_;
    Bit#(16) ipv4$totalLen;
  } IntAddUpdateVxlanGpeIpv4RspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_metadata_i2e$sink;
  } IntNoSinkRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) int_metadata$switch_id;
    Bit#(8) int_metadata$gpe_int_hdr_len8;
    Bit#(8) int_metadata$insert_cnt;
    Bit#(16) int_metadata$gpe_int_hdr_len;
    Bit#(16) int_metadata$insert_byte_cnt;
    Bit#(16) int_metadata$instruction_cnt;
  } IntResetRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_header$e;
  } IntSetEBitRspT;
  struct {
    PacketInstance pkt;
  } IntSetHeader0003I0RspT;
  struct {
    PacketInstance pkt;
    Bit#(24) int_q_occupancy_header$q_occupancy0;
    Bit#(7) int_q_occupancy_header$q_occupancy1;
  } IntSetHeader0003I1RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_switch_id_header$switch_id;
    Bit#(31) int_hop_latency_header$hop_latency;
  } IntSetHeader0003I10RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_switch_id_header$switch_id;
    Bit#(24) int_q_occupancy_header$q_occupancy0;
    Bit#(31) int_hop_latency_header$hop_latency;
    Bit#(7) int_q_occupancy_header$q_occupancy1;
  } IntSetHeader0003I11RspT;
  struct {
    PacketInstance pkt;
    Bit#(15) int_ingress_port_id_header$ingress_port_id_1;
    Bit#(16) int_ingress_port_id_header$ingress_port_id_0;
    Bit#(31) int_switch_id_header$switch_id;
  } IntSetHeader0003I12RspT;
  struct {
    PacketInstance pkt;
    Bit#(15) int_ingress_port_id_header$ingress_port_id_1;
    Bit#(24) int_q_occupancy_header$q_occupancy0;
    Bit#(16) int_ingress_port_id_header$ingress_port_id_0;
    Bit#(31) int_switch_id_header$switch_id;
    Bit#(7) int_q_occupancy_header$q_occupancy1;
  } IntSetHeader0003I13RspT;
  struct {
    PacketInstance pkt;
    Bit#(15) int_ingress_port_id_header$ingress_port_id_1;
    Bit#(16) int_ingress_port_id_header$ingress_port_id_0;
    Bit#(31) int_switch_id_header$switch_id;
    Bit#(31) int_hop_latency_header$hop_latency;
  } IntSetHeader0003I14RspT;
  struct {
    PacketInstance pkt;
    Bit#(24) int_q_occupancy_header$q_occupancy0;
    Bit#(31) int_switch_id_header$switch_id;
    Bit#(31) int_hop_latency_header$hop_latency;
    Bit#(15) int_ingress_port_id_header$ingress_port_id_1;
    Bit#(16) int_ingress_port_id_header$ingress_port_id_0;
    Bit#(7) int_q_occupancy_header$q_occupancy1;
  } IntSetHeader0003I15RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_hop_latency_header$hop_latency;
  } IntSetHeader0003I2RspT;
  struct {
    PacketInstance pkt;
    Bit#(24) int_q_occupancy_header$q_occupancy0;
    Bit#(31) int_hop_latency_header$hop_latency;
    Bit#(7) int_q_occupancy_header$q_occupancy1;
  } IntSetHeader0003I3RspT;
  struct {
    PacketInstance pkt;
    Bit#(15) int_ingress_port_id_header$ingress_port_id_1;
    Bit#(16) int_ingress_port_id_header$ingress_port_id_0;
  } IntSetHeader0003I4RspT;
  struct {
    PacketInstance pkt;
    Bit#(15) int_ingress_port_id_header$ingress_port_id_1;
    Bit#(24) int_q_occupancy_header$q_occupancy0;
    Bit#(16) int_ingress_port_id_header$ingress_port_id_0;
    Bit#(7) int_q_occupancy_header$q_occupancy1;
  } IntSetHeader0003I5RspT;
  struct {
    PacketInstance pkt;
    Bit#(15) int_ingress_port_id_header$ingress_port_id_1;
    Bit#(16) int_ingress_port_id_header$ingress_port_id_0;
    Bit#(31) int_hop_latency_header$hop_latency;
  } IntSetHeader0003I6RspT;
  struct {
    PacketInstance pkt;
    Bit#(15) int_ingress_port_id_header$ingress_port_id_1;
    Bit#(24) int_q_occupancy_header$q_occupancy0;
    Bit#(16) int_ingress_port_id_header$ingress_port_id_0;
    Bit#(31) int_hop_latency_header$hop_latency;
    Bit#(7) int_q_occupancy_header$q_occupancy1;
  } IntSetHeader0003I7RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_switch_id_header$switch_id;
  } IntSetHeader0003I8RspT;
  struct {
    PacketInstance pkt;
    Bit#(24) int_q_occupancy_header$q_occupancy0;
    Bit#(31) int_switch_id_header$switch_id;
    Bit#(7) int_q_occupancy_header$q_occupancy1;
  } IntSetHeader0003I9RspT;
  struct {
    PacketInstance pkt;
  } IntSetHeader0407I0RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_tx_utilization_header$egress_port_tx_utilization;
  } IntSetHeader0407I1RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_q_congestion_header$q_congestion;
    Bit#(31) int_ingress_tstamp_header$ingress_tstamp;
  } IntSetHeader0407I10RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_tx_utilization_header$egress_port_tx_utilization;
    Bit#(31) int_q_congestion_header$q_congestion;
    Bit#(31) int_ingress_tstamp_header$ingress_tstamp;
  } IntSetHeader0407I11RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_id_header$egress_port_id;
    Bit#(31) int_ingress_tstamp_header$ingress_tstamp;
  } IntSetHeader0407I12RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_tx_utilization_header$egress_port_tx_utilization;
    Bit#(31) int_egress_port_id_header$egress_port_id;
    Bit#(31) int_ingress_tstamp_header$ingress_tstamp;
  } IntSetHeader0407I13RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_q_congestion_header$q_congestion;
    Bit#(31) int_egress_port_id_header$egress_port_id;
    Bit#(31) int_ingress_tstamp_header$ingress_tstamp;
  } IntSetHeader0407I14RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_tx_utilization_header$egress_port_tx_utilization;
    Bit#(31) int_egress_port_id_header$egress_port_id;
    Bit#(31) int_q_congestion_header$q_congestion;
    Bit#(31) int_ingress_tstamp_header$ingress_tstamp;
  } IntSetHeader0407I15RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_q_congestion_header$q_congestion;
  } IntSetHeader0407I2RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_tx_utilization_header$egress_port_tx_utilization;
    Bit#(31) int_q_congestion_header$q_congestion;
  } IntSetHeader0407I3RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_id_header$egress_port_id;
  } IntSetHeader0407I4RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_tx_utilization_header$egress_port_tx_utilization;
    Bit#(31) int_egress_port_id_header$egress_port_id;
  } IntSetHeader0407I5RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_q_congestion_header$q_congestion;
    Bit#(31) int_egress_port_id_header$egress_port_id;
  } IntSetHeader0407I6RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_tx_utilization_header$egress_port_tx_utilization;
    Bit#(31) int_egress_port_id_header$egress_port_id;
    Bit#(31) int_q_congestion_header$q_congestion;
  } IntSetHeader0407I7RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_ingress_tstamp_header$ingress_tstamp;
  } IntSetHeader0407I8RspT;
  struct {
    PacketInstance pkt;
    Bit#(31) int_egress_port_tx_utilization_header$egress_port_tx_utilization;
    Bit#(31) int_ingress_tstamp_header$ingress_tstamp;
  } IntSetHeader0407I9RspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_switch_id_header$bos;
  } IntSetHeader0BosRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_ingress_port_id_header$bos;
  } IntSetHeader1BosRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_hop_latency_header$bos;
  } IntSetHeader2BosRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_q_occupancy_header$bos;
  } IntSetHeader3BosRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_ingress_tstamp_header$bos;
  } IntSetHeader4BosRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_egress_port_id_header$bos;
  } IntSetHeader5BosRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_q_congestion_header$bos;
  } IntSetHeader6BosRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_egress_port_tx_utilization_header$bos;
  } IntSetHeader7BosRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_metadata_i2e$source;
  } IntSetNoSrcRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) int_metadata_i2e$source;
  } IntSetSrcRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) i2e_metadata$mirror_session_id;
    Bit#(1) int_metadata_i2e$sink;
  } IntSinkGpeRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) vxlan_gpe$next_proto;
  } IntSinkUpdateVxlanGpeV4RspT;
  struct {
    PacketInstance pkt;
    Bit#(8) int_metadata$gpe_int_hdr_len8;
    Bit#(16) int_header$rsvd2;
    Bit#(5) int_header$ins_cnt;
    Bit#(4) int_header$instruction_mask_0407;
    Bit#(8) int_header$total_hop_cnt;
    Bit#(4) int_header$instruction_mask_1215;
    Bit#(5) int_header$rsvd1;
    Bit#(1) int_header$e;
    Bit#(4) int_header$instruction_mask_0811;
    Bit#(32) int_metadata$switch_id;
    Bit#(2) int_header$rep;
    Bit#(2) int_header$ver;
    Bit#(8) int_header$max_hop_cnt;
    Bit#(4) int_header$instruction_mask_0003;
    Bit#(8) int_metadata$insert_cnt;
    Bit#(1) int_header$c;
    Bit#(16) int_metadata$insert_byte_cnt;
  } IntSrcRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) int_metadata$switch_id;
    Bit#(8) int_metadata$gpe_int_hdr_len8;
  } IntTransitRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) int_header$total_hop_cnt;
  } IntUpdateTotalHopCntRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) vxlan_gpe_int_header$len;
    Bit#(16) udp$length_;
    Bit#(16) ipv4$totalLen;
  } IntUpdateVxlanGpeIpv4RspT;
  struct {
    PacketInstance pkt;
    Bit#(1) security_metadata$ipsg_check_fail;
  } IpsgMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) gre$S;
    Bit#(16) ipv4$identification;
    Bit#(1) gre$s;
    Bit#(4) ipv4$version;
    Bit#(4) ipv4$ihl;
    Bit#(16) gre$proto;
    Bit#(8) ipv4$ttl;
    Bit#(3) gre$ver;
    Bit#(32) erspan_t3_header$timestamp;
    Bit#(1) gre$C;
    Bit#(3) gre$recurse;
    Bit#(10) erspan_t3_header$span_id;
    Bit#(1) gre$K;
    Bit#(4) erspan_t3_header$version;
    Bit#(5) gre$flags;
    Bit#(32) erspan_t3_header$sgt_other;
    Bit#(8) ipv4$protocol;
    Bit#(1) gre$R;
  } Ipv4ErspanT3RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(24) genv$vni;
    Bit#(16) ipv4$identification;
    Bit#(16) udp$checksum;
    Bit#(4) ipv4$version;
    Bit#(4) ipv4$ihl;
    Bit#(6) genv$optLen;
    Bit#(8) ipv4$ttl;
    Bit#(1) genv$oam;
    Bit#(8) genv$reserved2;
    Bit#(1) genv$critical;
    Bit#(16) udp$srcPort;
    Bit#(16) genv$protoType;
    Bit#(2) genv$ver;
    Bit#(16) udp$dstPort;
    Bit#(16) ethernet$etherType;
    Bit#(8) ipv4$protocol;
    Bit#(6) genv$reserved;
  } Ipv4GenvRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ipv4$protocol;
    Bit#(4) ipv4$ihl;
    Bit#(16) gre$proto;
    Bit#(8) ipv4$ttl;
    Bit#(16) ipv4$identification;
    Bit#(16) ethernet$etherType;
    Bit#(4) ipv4$version;
  } Ipv4GreRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ipv4$protocol;
    Bit#(4) ipv4$ihl;
    Bit#(8) ipv4$ttl;
    Bit#(16) ipv4$identification;
    Bit#(16) ethernet$etherType;
    Bit#(4) ipv4$version;
  } Ipv4IpRewriteRspT;
  struct {
    PacketInstance pkt;
  } Ipv4MtuCheckRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ipv4$ttl;
  } Ipv4MulticastRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) gre$s;
    Bit#(16) ipv4$identification;
    Bit#(1) gre$R;
    Bit#(8) nvgre$flow_id;
    Bit#(4) ipv4$ihl;
    Bit#(16) gre$proto;
    Bit#(8) ipv4$ttl;
    Bit#(3) gre$ver;
    Bit#(1) gre$S;
    Bit#(1) gre$C;
    Bit#(3) gre$recurse;
    Bit#(24) nvgre$tni;
    Bit#(1) gre$K;
    Bit#(5) gre$flags;
    Bit#(16) ethernet$etherType;
    Bit#(8) ipv4$protocol;
    Bit#(4) ipv4$version;
  } Ipv4NvgreRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) ipv4_metadata$lkp_ipv4_da;
    Bit#(32) ipv4_metadata$lkp_ipv4_sa;
    Bit#(16) l3_metadata$lkp_l4_dport;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(16) l3_metadata$lkp_l4_sport;
    Bit#(8) l3_metadata$lkp_ip_proto;
    Bit#(48) l2_metadata$lkp_mac_da;
  } Ipv4OverFabricRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) l3_metadata$lkp_ip_ttl;
    Bit#(32) ipv4_metadata$lkp_ipv4_da;
    Bit#(32) ipv4_metadata$lkp_ipv4_sa;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(16) l3_metadata$lkp_l4_dport;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(16) l3_metadata$lkp_l4_sport;
    Bit#(8) l3_metadata$lkp_ip_proto;
    Bit#(48) l2_metadata$lkp_mac_da;
  } Ipv4TunnelLookupMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ipv4$ttl;
    Bit#(48) ethernet$dstAddr;
  } Ipv4UnicastRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$urpf_bd_group;
    Bit#(1) l3_metadata$urpf_hit;
    Bit#(2) l3_metadata$urpf_mode;
  } Ipv4UrpfHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ipv4$identification;
    Bit#(16) udp$checksum;
    Bit#(None) vxlan$vni;
    Bit#(4) ipv4$ihl;
    Bit#(None) vxlan$flags;
    Bit#(8) ipv4$ttl;
    Bit#(8) ipv4$protocol;
    Bit#(None) vxlan$reserved2;
    Bit#(16) udp$srcPort;
    Bit#(None) vxlan$reserved;
    Bit#(16) udp$dstPort;
    Bit#(16) ethernet$etherType;
    Bit#(4) ipv4$version;
  } Ipv4VxlanRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ipv6$version;
    Bit#(1) gre$S;
    Bit#(8) ipv6$trafficClass;
    Bit#(1) gre$s;
    Bit#(8) ipv6$hopLimit;
    Bit#(20) ipv6$flowLabel;
    Bit#(16) gre$proto;
    Bit#(3) gre$ver;
    Bit#(32) erspan_t3_header$timestamp;
    Bit#(1) gre$C;
    Bit#(3) gre$recurse;
    Bit#(8) ipv6$nextHdr;
    Bit#(10) erspan_t3_header$span_id;
    Bit#(1) gre$K;
    Bit#(4) erspan_t3_header$version;
    Bit#(5) gre$flags;
    Bit#(32) erspan_t3_header$sgt_other;
    Bit#(1) gre$R;
  } Ipv6ErspanT3RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(24) genv$vni;
    Bit#(8) ipv6$trafficClass;
    Bit#(16) udp$checksum;
    Bit#(4) ipv6$version;
    Bit#(6) genv$optLen;
    Bit#(8) ipv6$nextHdr;
    Bit#(1) genv$oam;
    Bit#(8) genv$reserved2;
    Bit#(16) ethernet$etherType;
    Bit#(1) genv$critical;
    Bit#(16) udp$srcPort;
    Bit#(20) ipv6$flowLabel;
    Bit#(16) genv$protoType;
    Bit#(2) genv$ver;
    Bit#(16) udp$dstPort;
    Bit#(8) ipv6$hopLimit;
    Bit#(6) genv$reserved;
  } Ipv6GenvRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ipv6$version;
    Bit#(20) ipv6$flowLabel;
    Bit#(16) gre$proto;
    Bit#(8) ipv6$hopLimit;
    Bit#(8) ipv6$trafficClass;
    Bit#(8) ipv6$nextHdr;
    Bit#(16) ethernet$etherType;
  } Ipv6GreRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ipv6$version;
    Bit#(16) ipv6$payloadLen;
    Bit#(20) ipv6$flowLabel;
    Bit#(8) ipv6$hopLimit;
    Bit#(8) ipv6$trafficClass;
    Bit#(8) ipv6$nextHdr;
    Bit#(16) ethernet$etherType;
  } Ipv6IpRewriteRspT;
  struct {
    PacketInstance pkt;
  } Ipv6MtuCheckRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ipv6$hopLimit;
  } Ipv6MulticastRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ipv6$version;
    Bit#(1) gre$s;
    Bit#(1) gre$R;
    Bit#(8) nvgre$flow_id;
    Bit#(16) gre$proto;
    Bit#(3) gre$ver;
    Bit#(1) gre$S;
    Bit#(16) ethernet$etherType;
    Bit#(1) gre$C;
    Bit#(3) gre$recurse;
    Bit#(24) nvgre$tni;
    Bit#(8) ipv6$nextHdr;
    Bit#(20) ipv6$flowLabel;
    Bit#(1) gre$K;
    Bit#(8) ipv6$trafficClass;
    Bit#(5) gre$flags;
    Bit#(8) ipv6$hopLimit;
  } Ipv6NvgreRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(128) ipv6_metadata$lkp_ipv6_sa;
    Bit#(128) ipv6_metadata$lkp_ipv6_da;
    Bit#(16) l3_metadata$lkp_l4_sport;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(16) l3_metadata$lkp_l4_dport;
    Bit#(8) l3_metadata$lkp_ip_proto;
    Bit#(48) l2_metadata$lkp_mac_da;
  } Ipv6OverFabricRspT;
  struct {
    PacketInstance pkt;
    Bit#(128) ipv6_metadata$lkp_ipv6_sa;
    Bit#(128) ipv6_metadata$lkp_ipv6_da;
    Bit#(16) l3_metadata$lkp_l4_sport;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(8) l3_metadata$lkp_ip_ttl;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(16) l3_metadata$lkp_l4_dport;
    Bit#(8) l3_metadata$lkp_ip_proto;
    Bit#(48) l2_metadata$lkp_mac_da;
  } Ipv6TunnelLookupMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ipv6$hopLimit;
    Bit#(48) ethernet$dstAddr;
  } Ipv6UnicastRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$urpf_bd_group;
    Bit#(1) l3_metadata$urpf_hit;
    Bit#(2) l3_metadata$urpf_mode;
  } Ipv6UrpfHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ipv6$version;
    Bit#(16) udp$checksum;
    Bit#(None) vxlan$vni;
    Bit#(None) vxlan$flags;
    Bit#(8) ipv6$nextHdr;
    Bit#(None) vxlan$reserved2;
    Bit#(16) udp$srcPort;
    Bit#(20) ipv6$flowLabel;
    Bit#(None) vxlan$reserved;
    Bit#(8) ipv6$hopLimit;
    Bit#(8) ipv6$trafficClass;
    Bit#(16) udp$dstPort;
    Bit#(16) ethernet$etherType;
  } Ipv6VxlanRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ingress_metadata$drop_reason;
    Bit#(1) ingress_metadata$drop_flag;
  } MalformedOuterEthernetPacketRspT;
  struct {
    PacketInstance pkt;
  } MeterDenyRspT;
  struct {
    PacketInstance pkt;
  } MeterPermitRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } MplsEthernetPush1RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } MplsEthernetPush2RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } MplsEthernetPush3RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } MplsIpPush1RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } MplsIpPush2RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } MplsIpPush3RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$dstAddr;
    Bit#(8) mpls0$ttl;
  } MplsRewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$l3_mtu_check;
  } MtuMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) multicast_metadata$mcast_bridge_hit;
    Bit#(16) multicast_metadata$multicast_bridge_mc_index;
  } MulticastBridgeSGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) multicast_metadata$mcast_bridge_hit;
    Bit#(16) multicast_metadata$multicast_bridge_mc_index;
  } MulticastBridgeStarGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) multicast_metadata$mcast_route_hit;
    Bit#(16) multicast_metadata$multicast_route_mc_index;
    Bit#(2) multicast_metadata$mcast_mode;
  } MulticastRouteBidirStarGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) multicast_metadata$mcast_route_hit;
    Bit#(16) multicast_metadata$multicast_route_mc_index;
    Bit#(2) multicast_metadata$mcast_mode;
  } MulticastRouteSGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) multicast_metadata$mcast_route_hit;
    Bit#(16) multicast_metadata$multicast_route_mc_index;
    Bit#(2) multicast_metadata$mcast_mode;
  } MulticastRouteSmStarGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$l3_copy;
  } MulticastRouteStarGMissRspT;
  struct {
    PacketInstance pkt;
  } NegativeMirrorRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(16) l2_metadata$lkp_mac_type;
    Bit#(48) l2_metadata$lkp_mac_da;
  } NonIpOverFabricRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(48) l2_metadata$lkp_mac_da;
  } NonIpTunnelLookupMissRspT;
  struct {
    PacketInstance pkt;
  } NopRspT;
  struct {
    PacketInstance pkt;
  } OnMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } OuterMulticastBridgeSGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } OuterMulticastBridgeStarGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(1) multicast_metadata$outer_mcast_route_hit;
    Bit#(2) multicast_metadata$outer_mcast_mode;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } OuterMulticastRouteBidirStarGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(1) multicast_metadata$outer_mcast_route_hit;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } OuterMulticastRouteSGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(1) multicast_metadata$outer_mcast_route_hit;
    Bit#(2) multicast_metadata$outer_mcast_mode;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } OuterMulticastRouteSmStarGHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) multicast_metadata$replica;
    Bit#(1) multicast_metadata$inner_replica;
    Bit#(4) tunnel_metadata$egress_header_count;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
    Bit#(16) egress_metadata$bd;
    Bit#(14) tunnel_metadata$tunnel_index;
    Bit#(1) egress_metadata$routed;
  } OuterReplicaFromRidRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$rmac_hit;
  } OuterRmacHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l2_metadata$port_vlan_mapping_miss;
  } PortVlanMappingMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) acl_metadata$racl_deny;
    Bit#(1) acl_metadata$acl_copy;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(14) acl_metadata$acl_stats_index;
  } RaclDenyRspT;
  struct {
    PacketInstance pkt;
    Bit#(14) acl_metadata$acl_stats_index;
    Bit#(1) acl_metadata$acl_copy;
    Bit#(16) fabric_metadata$reason_code;
  } RaclPermitRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) acl_metadata$racl_nexthop;
    Bit#(1) acl_metadata$acl_copy;
    Bit#(14) acl_metadata$acl_stats_index;
    Bit#(1) acl_metadata$racl_redirect;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(1) acl_metadata$racl_nexthop_type;
  } RaclRedirectEcmpRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) acl_metadata$racl_nexthop;
    Bit#(1) acl_metadata$acl_copy;
    Bit#(14) acl_metadata$acl_stats_index;
    Bit#(1) acl_metadata$racl_redirect;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(1) acl_metadata$racl_nexthop_type;
  } RaclRedirectNexthopRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) fabric_metadata$reason_code;
  } RedirectToCpuRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } RemoveVlanDoubleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ethernet$etherType;
  } RemoveVlanSingleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$dstAddr;
  } RewriteIpv4MulticastRspT;
  struct {
    PacketInstance pkt;
  } RewriteIpv6MulticastRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
  } RewriteSmacRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$dstAddr;
  } RewriteTunnelDmacRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) ipv4$dstAddr;
  } RewriteTunnelIpv4DstRspT;
  struct {
    PacketInstance pkt;
    Bit#(32) ipv4$srcAddr;
  } RewriteTunnelIpv4SrcRspT;
  struct {
    PacketInstance pkt;
    Bit#(128) ipv6$dstAddr;
  } RewriteTunnelIpv6DstRspT;
  struct {
    PacketInstance pkt;
    Bit#(128) ipv6$srcAddr;
  } RewriteTunnelIpv6SrcRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) ethernet$srcAddr;
  } RewriteTunnelSmacRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$rmac_hit;
  } RmacHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$rmac_hit;
  } RmacMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(1) nexthop_metadata$nexthop_type;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetAclRedirectActionRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } SetBdFloodMcIndexRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) multicast_metadata$ipv4_mcast_key;
    Bit#(10) l3_metadata$rmac_group;
    Bit#(1) multicast_metadata$igmp_snooping_enabled;
    Bit#(16) multicast_metadata$bd_mrpf_group;
    Bit#(1) multicast_metadata$ipv4_multicast_enabled;
    Bit#(1) multicast_metadata$mld_snooping_enabled;
    Bit#(16) acl_metadata$bd_label;
    Bit#(10) l2_metadata$stp_group;
    Bit#(16) l3_metadata$vrf;
    Bit#(2) ipv6_metadata$ipv6_urpf_mode;
    Bit#(1) ipv6_metadata$ipv6_unicast_enabled;
    Bit#(1) l2_metadata$learning_enabled;
    Bit#(16) ingress_metadata$outer_bd;
    Bit#(16) multicast_metadata$ipv6_mcast_key;
    Bit#(16) ingress_metadata$bd;
    Bit#(1) multicast_metadata$ipv4_mcast_key_type;
    Bit#(1) multicast_metadata$ipv6_mcast_key_type;
    Bit#(2) ipv4_metadata$ipv4_urpf_mode;
    Bit#(1) multicast_metadata$ipv6_multicast_enabled;
    Bit#(16) l2_metadata$bd_stats_idx;
    Bit#(1) ipv4_metadata$ipv4_unicast_enabled;
  } SetBdPropertiesRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$bd_stats_idx;
  } SetBroadcastRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) intrinsic_metadata$deflect_on_drop;
    Bit#(32) i2e_metadata$ingress_tstamp;
    Bit#(9) ingress_metadata$ingress_port;
    Bit#(9) standard_metadata$egress_spec;
    Bit#(16) l2_metadata$same_if_check;
  } SetConfigParametersRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$routed;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) ingress_metadata$egress_ifindex;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(9) standard_metadata$egress_spec;
  } SetCpuRedirectActionRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetEcmpNexthopDetailsRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetEcmpNexthopDetailsForPostRoutedFloodRspT;
  struct {
    PacketInstance pkt;
    Bit#(9) egress_metadata$smac_idx;
  } SetEgressBdPropertiesRspT;
  struct {
    PacketInstance pkt;
  } SetEgressFilterDropRspT;
  struct {
    PacketInstance pkt;
    Bit#(12) vlan_tag_1$vid;
    Bit#(12) vlan_tag_0$vid;
    Bit#(16) vlan_tag_0$etherType;
    Bit#(16) vlan_tag_1$etherType;
    Bit#(16) ethernet$etherType;
  } SetEgressPacketVlanDoubleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(12) vlan_tag_0$vid;
    Bit#(16) vlan_tag_0$etherType;
    Bit#(16) ethernet$etherType;
  } SetEgressPacketVlanTaggedRspT;
  struct {
    PacketInstance pkt;
  } SetEgressPacketVlanUntaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(24) tunnel_metadata$vnid;
  } SetEgressTunnelVniRspT;
  struct {
    PacketInstance pkt;
    Bit#(9) standard_metadata$egress_spec;
  } SetFabricLagPortRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) multicast_metadata$mcast_grp;
  } SetFabricMulticastRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(1) nexthop_metadata$nexthop_type;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(1) l3_metadata$routed;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) fabric_metadata$reason_code;
  } SetFibRedirectActionRspT;
  struct {
    PacketInstance pkt;
    Bit#(2) ingress_metadata$port_type;
    Bit#(16) ingress_metadata$ifindex;
  } SetIfindexRspT;
  struct {
    PacketInstance pkt;
  } SetIngressIfindexPropertiesRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) acl_metadata$if_label;
  } SetIngressPortPropertiesRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(1) nexthop_metadata$nexthop_type;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetL2RedirectActionRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$outer_bd;
    Bit#(16) egress_metadata$bd;
    Bit#(1) egress_metadata$routed;
  } SetL2RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$outer_bd;
    Bit#(16) egress_metadata$bd;
    Bit#(14) tunnel_metadata$tunnel_index;
    Bit#(1) egress_metadata$routed;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
  } SetL2RewriteWithTunnelRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$outer_bd;
    Bit#(16) egress_metadata$bd;
    Bit#(48) egress_metadata$mac_da;
    Bit#(1) egress_metadata$routed;
    Bit#(8) l3_metadata$mtu_index;
  } SetL3RewriteRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$outer_bd;
    Bit#(14) tunnel_metadata$tunnel_index;
    Bit#(48) egress_metadata$mac_da;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
    Bit#(16) egress_metadata$bd;
    Bit#(1) egress_metadata$routed;
  } SetL3RewriteWithTunnelRspT;
  struct {
    PacketInstance pkt;
  } SetLagMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(9) standard_metadata$egress_spec;
  } SetLagPortRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) fabric_metadata$dst_port;
  } SetLagRemotePortRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ingress_metadata$drop_reason;
    Bit#(1) ingress_metadata$drop_flag;
  } SetMalformedOuterIpv4PacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ingress_metadata$drop_reason;
    Bit#(1) ingress_metadata$drop_flag;
  } SetMalformedOuterIpv6PacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ingress_metadata$drop_reason;
    Bit#(1) ingress_metadata$drop_flag;
  } SetMalformedPacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$bd;
  } SetMirrorBdRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
  } SetMirrorNhopRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$bd;
    Bit#(14) tunnel_metadata$tunnel_index;
    Bit#(4) tunnel_metadata$egress_header_count;
    Bit#(1) egress_metadata$routed;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
  } SetMplsPushRewriteL2RspT;
  struct {
    PacketInstance pkt;
    Bit#(14) tunnel_metadata$tunnel_index;
    Bit#(1) egress_metadata$routed;
    Bit#(48) egress_metadata$mac_da;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
    Bit#(16) egress_metadata$bd;
    Bit#(4) tunnel_metadata$egress_header_count;
  } SetMplsPushRewriteL3RspT;
  struct {
    PacketInstance pkt;
    Bit#(9) tunnel_metadata$tunnel_smac_index;
    Bit#(3) mpls0$exp;
    Bit#(8) mpls0$ttl;
    Bit#(1) mpls0$bos;
    Bit#(14) tunnel_metadata$tunnel_dmac_index;
    Bit#(20) mpls0$label;
  } SetMplsRewritePush1RspT;
  struct {
    PacketInstance pkt;
    Bit#(8) mpls1$ttl;
    Bit#(9) tunnel_metadata$tunnel_smac_index;
    Bit#(3) mpls1$exp;
    Bit#(3) mpls0$exp;
    Bit#(8) mpls0$ttl;
    Bit#(20) mpls1$label;
    Bit#(1) mpls0$bos;
    Bit#(1) mpls1$bos;
    Bit#(14) tunnel_metadata$tunnel_dmac_index;
    Bit#(20) mpls0$label;
  } SetMplsRewritePush2RspT;
  struct {
    PacketInstance pkt;
    Bit#(8) mpls1$ttl;
    Bit#(3) mpls1$exp;
    Bit#(1) mpls2$bos;
    Bit#(9) tunnel_metadata$tunnel_smac_index;
    Bit#(20) mpls1$label;
    Bit#(1) mpls0$bos;
    Bit#(3) mpls2$exp;
    Bit#(8) mpls2$ttl;
    Bit#(3) mpls0$exp;
    Bit#(14) tunnel_metadata$tunnel_dmac_index;
    Bit#(8) mpls0$ttl;
    Bit#(20) mpls2$label;
    Bit#(1) mpls1$bos;
    Bit#(20) mpls0$label;
  } SetMplsRewritePush3RspT;
  struct {
    PacketInstance pkt;
    Bit#(14) tunnel_metadata$tunnel_index;
    Bit#(1) egress_metadata$routed;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
    Bit#(16) egress_metadata$bd;
    Bit#(4) tunnel_metadata$egress_header_count;
    Bit#(20) mpls0$label;
  } SetMplsSwapPushRewriteL2RspT;
  struct {
    PacketInstance pkt;
    Bit#(14) tunnel_metadata$tunnel_index;
    Bit#(4) tunnel_metadata$egress_header_count;
    Bit#(48) egress_metadata$mac_da;
    Bit#(5) tunnel_metadata$egress_tunnel_type;
    Bit#(16) egress_metadata$bd;
    Bit#(1) egress_metadata$routed;
    Bit#(20) mpls0$label;
  } SetMplsSwapPushRewriteL3RspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$bd_stats_idx;
  } SetMulticastRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(1) ipv6_metadata$ipv6_src_is_link_local;
    Bit#(16) l2_metadata$bd_stats_idx;
  } SetMulticastAndIpv6SrcIsLinkLocalRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetMulticastBridgeActionRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ingress_metadata$drop_reason;
    Bit#(1) ingress_metadata$drop_flag;
  } SetMulticastDropRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetMulticastFloodRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$routed;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(16) l3_metadata$same_bd_check;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetMulticastRouteActionRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetNexthopDetailsRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) fabric_metadata$dst_device;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(16) ingress_metadata$egress_ifindex;
  } SetNexthopDetailsForPostRoutedFloodRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(1) nexthop_metadata$nexthop_type;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(16) ingress_metadata$egress_ifindex;
    Bit#(1) l3_metadata$routed;
    Bit#(8) fabric_metadata$dst_device;
  } SetRaclRedirectActionRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) egress_metadata$routed;
  } SetReplicaCopyBridgedRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) meter_metadata$meter_index;
  } SetStormControlMeterRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$stp_state;
  } SetStpStateRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) egress_metadata$outer_bd;
    Bit#(9) tunnel_metadata$tunnel_src_index;
    Bit#(14) tunnel_metadata$tunnel_dst_index;
    Bit#(14) tunnel_metadata$tunnel_dmac_index;
    Bit#(9) tunnel_metadata$tunnel_smac_index;
  } SetTunnelRewriteDetailsRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) tunnel_metadata$tunnel_terminate;
  } SetTunnelTerminationFlagRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(24) tunnel_metadata$tunnel_vni;
  } SetTunnelVniAndTerminationFlagRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
  } SetUnicastRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(1) ipv6_metadata$ipv6_src_is_link_local;
  } SetUnicastAndIpv6SrcIsLinkLocalRspT;
  struct {
    PacketInstance pkt;
    Bit#(20) tunnel_metadata$mpls_label;
    Bit#(3) tunnel_metadata$mpls_exp;
  } SetValidMplsLabel1RspT;
  struct {
    PacketInstance pkt;
    Bit#(20) tunnel_metadata$mpls_label;
    Bit#(3) tunnel_metadata$mpls_exp;
  } SetValidMplsLabel2RspT;
  struct {
    PacketInstance pkt;
    Bit#(20) tunnel_metadata$mpls_label;
    Bit#(3) tunnel_metadata$mpls_exp;
  } SetValidMplsLabel3RspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterBroadcastPacketDoubleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterBroadcastPacketQinqTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterBroadcastPacketSingleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterBroadcastPacketUntaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(4) l3_metadata$lkp_ip_version;
  } SetValidOuterIpv4PacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(4) l3_metadata$lkp_ip_version;
  } SetValidOuterIpv6PacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterMulticastPacketDoubleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterMulticastPacketQinqTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterMulticastPacketSingleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterMulticastPacketUntaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterUnicastPacketDoubleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterUnicastPacketQinqTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterUnicastPacketSingleTaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(3) l2_metadata$lkp_pkt_type;
    Bit#(16) l2_metadata$lkp_mac_type;
  } SetValidOuterUnicastPacketUntaggedRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) fabric_metadata$reason_code;
    Bit#(16) i2e_metadata$mirror_session_id;
  } SflowIngPktToCpuRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) sflow_metadata$sflow_session_id;
  } SflowIngSessionEnableRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) fabric_header_sflow$sflow_session_id;
  } SflowPktToCpuRspT;
  struct {
    PacketInstance pkt;
  } SmacHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l2_metadata$l2_src_miss;
  } SmacMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) ingress_metadata$ifindex;
  } SrcVtepHitRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) fabric_metadata$fabric_header_present;
    Bit#(16) intrinsic_metadata$mcast_grp;
  } SwitchFabricMulticastPacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) fabric_metadata$fabric_header_present;
    Bit#(16) fabric_metadata$dst_port;
    Bit#(8) fabric_metadata$dst_device;
  } SwitchFabricUnicastPacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) egress_metadata$bypass;
    Bit#(9) standard_metadata$egress_spec;
    Bit#(16) ethernet$etherType;
  } TerminateCpuPacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(5) tunnel_metadata$ingress_tunnel_type;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) l2_metadata$lkp_mac_type;
    Bit#(16) ingress_metadata$bd;
  } TerminateEomplsRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(5) tunnel_metadata$ingress_tunnel_type;
    Bit#(16) intrinsic_metadata$mcast_grp;
    Bit#(1) l3_metadata$routed;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) ethernet$etherType;
    Bit#(1) l3_metadata$outer_routed;
  } TerminateFabricMulticastPacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$nexthop_index;
    Bit#(5) tunnel_metadata$ingress_tunnel_type;
    Bit#(9) standard_metadata$egress_spec;
    Bit#(1) l3_metadata$routed;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) ethernet$etherType;
    Bit#(1) l3_metadata$outer_routed;
  } TerminateFabricUnicastPacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(5) tunnel_metadata$ingress_tunnel_type;
    Bit#(16) l2_metadata$lkp_mac_type;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) l3_metadata$vrf;
    Bit#(4) l3_metadata$lkp_ip_version;
    Bit#(48) l2_metadata$lkp_mac_da;
  } TerminateIpv4OverMplsRspT;
  struct {
    PacketInstance pkt;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(5) tunnel_metadata$ingress_tunnel_type;
    Bit#(16) l2_metadata$lkp_mac_type;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) l3_metadata$vrf;
    Bit#(4) l3_metadata$lkp_ip_version;
    Bit#(48) l2_metadata$lkp_mac_da;
  } TerminateIpv6OverMplsRspT;
  struct {
    PacketInstance pkt;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(48) l2_metadata$lkp_mac_da;
    Bit#(16) ingress_metadata$egress_ifindex;
  } TerminatePwRspT;
  struct {
    PacketInstance pkt;
    Bit#(10) l3_metadata$rmac_group;
    Bit#(1) multicast_metadata$igmp_snooping_enabled;
    Bit#(16) multicast_metadata$bd_mrpf_group;
    Bit#(1) multicast_metadata$ipv4_multicast_enabled;
    Bit#(16) l2_metadata$lkp_mac_type;
    Bit#(16) acl_metadata$bd_label;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(16) l3_metadata$vrf;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(4) l3_metadata$lkp_ip_version;
    Bit#(8) qos_metadata$outer_dscp;
    Bit#(16) ingress_metadata$bd;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(2) ipv4_metadata$ipv4_urpf_mode;
    Bit#(16) l2_metadata$bd_stats_idx;
    Bit#(1) ipv4_metadata$ipv4_unicast_enabled;
  } TerminateTunnelInnerEthernetIpv4RspT;
  struct {
    PacketInstance pkt;
    Bit#(10) l3_metadata$rmac_group;
    Bit#(16) multicast_metadata$bd_mrpf_group;
    Bit#(16) l2_metadata$lkp_mac_type;
    Bit#(16) acl_metadata$bd_label;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(16) l3_metadata$vrf;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(1) ipv6_metadata$ipv6_unicast_enabled;
    Bit#(2) ipv6_metadata$ipv6_urpf_mode;
    Bit#(8) qos_metadata$outer_dscp;
    Bit#(16) ingress_metadata$bd;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(1) multicast_metadata$ipv6_multicast_enabled;
    Bit#(16) l2_metadata$bd_stats_idx;
    Bit#(4) l3_metadata$lkp_ip_version;
    Bit#(1) multicast_metadata$mld_snooping_enabled;
  } TerminateTunnelInnerEthernetIpv6RspT;
  struct {
    PacketInstance pkt;
    Bit#(10) l3_metadata$rmac_group;
    Bit#(2) ipv4_metadata$ipv4_urpf_mode;
    Bit#(16) multicast_metadata$bd_mrpf_group;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(16) l3_metadata$vrf;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(1) multicast_metadata$ipv4_multicast_enabled;
    Bit#(8) qos_metadata$outer_dscp;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(1) ipv4_metadata$ipv4_unicast_enabled;
    Bit#(4) l3_metadata$lkp_ip_version;
    Bit#(48) l2_metadata$lkp_mac_da;
  } TerminateTunnelInnerIpv4RspT;
  struct {
    PacketInstance pkt;
    Bit#(10) l3_metadata$rmac_group;
    Bit#(8) qos_metadata$outer_dscp;
    Bit#(16) multicast_metadata$bd_mrpf_group;
    Bit#(48) l2_metadata$lkp_mac_sa;
    Bit#(8) l3_metadata$lkp_ip_tc;
    Bit#(16) l3_metadata$vrf;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(1) ipv6_metadata$ipv6_unicast_enabled;
    Bit#(128) ipv6_metadata$lkp_ipv6_sa;
    Bit#(2) ipv6_metadata$ipv6_urpf_mode;
    Bit#(128) ipv6_metadata$lkp_ipv6_da;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(1) multicast_metadata$ipv6_multicast_enabled;
    Bit#(4) l3_metadata$lkp_ip_version;
    Bit#(48) l2_metadata$lkp_mac_da;
  } TerminateTunnelInnerIpv6RspT;
  struct {
    PacketInstance pkt;
    Bit#(2) l3_metadata$lkp_ip_type;
    Bit#(16) ingress_metadata$bd;
    Bit#(16) l2_metadata$lkp_mac_type;
    Bit#(16) acl_metadata$bd_label;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) l2_metadata$bd_stats_idx;
  } TerminateTunnelInnerNonIpRspT;
  struct {
    PacketInstance pkt;
    Bit#(5) tunnel_metadata$ingress_tunnel_type;
    Bit#(1) tunnel_metadata$tunnel_terminate;
    Bit#(16) l2_metadata$lkp_mac_type;
    Bit#(16) ingress_metadata$bd;
  } TerminateVplsRspT;
  struct {
    PacketInstance pkt;
  } TunnelLookupMissRspT;
  struct {
    PacketInstance pkt;
  } TunnelMtuCheckRspT;
  struct {
    PacketInstance pkt;
    Bit#(16) l3_metadata$l3_mtu_check;
  } TunnelMtuMissRspT;
  struct {
    PacketInstance pkt;
  } UpdateIngressBdStatsRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$urpf_check_fail;
  } UrpfBdMissRspT;
  struct {
    PacketInstance pkt;
    Bit#(1) l3_metadata$urpf_check_fail;
  } UrpfMissRspT;
} BBResponse deriving (Bits, Eq, FShow);

// ====== ACL_DENY ======

interface AclDeny;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkAclDeny  (AclDeny);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) acl_metadata$acl_deny <- mkReg(0);
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(16)) meter_metadata$meter_index <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_copy <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule acl_deny_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged AclDenyReqT {pkt: .pkt, runtime_acl_copy_reason: .runtime_acl_copy_reason, runtime_acl_copy: .runtime_acl_copy, runtime_acl_meter_index: .runtime_acl_meter_index, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        acl_metadata$acl_deny <= 'h1;
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        meter_metadata$meter_index <= runtime_acl_meter_index;
        acl_metadata$acl_copy <= runtime_acl_copy;
        fabric_metadata$reason_code <= runtime_acl_copy_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule acl_deny_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged AclDenyRspT {pkt: pkt, acl_metadata$acl_deny: acl_metadata$acl_deny, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index, meter_metadata$meter_index: meter_metadata$meter_index, fabric_metadata$reason_code: fabric_metadata$reason_code, acl_metadata$acl_copy: acl_metadata$acl_copy};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== ACL_MIRROR ======

interface AclMirror;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkAclMirror  (AclMirror);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) i2e_metadata$mirror_session_id <- mkReg(0);
  Reg#(Bit#(32)) i2e_metadata$ingress_tstamp <- mkReg(0);
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(16)) meter_metadata$meter_index <- mkReg(0);
  rule acl_mirror_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged AclMirrorReqT {pkt: .pkt, intrinsic_metadata$ingress_global_tstamp: .intrinsic_metadata$ingress_global_tstamp, runtime_session_id: .runtime_session_id, runtime_acl_meter_index: .runtime_acl_meter_index, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        i2e_metadata$mirror_session_id <= runtime_session_id;
        i2e_metadata$ingress_tstamp <= intrinsic_metadata$ingress_global_tstamp;
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        meter_metadata$meter_index <= runtime_acl_meter_index;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule acl_mirror_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged AclMirrorRspT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index, meter_metadata$meter_index: meter_metadata$meter_index, i2e_metadata$mirror_session_id: i2e_metadata$mirror_session_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== ACL_PERMIT ======

interface AclPermit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkAclPermit  (AclPermit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(16)) meter_metadata$meter_index <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_copy <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule acl_permit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged AclPermitReqT {pkt: .pkt, runtime_acl_copy_reason: .runtime_acl_copy_reason, runtime_acl_copy: .runtime_acl_copy, runtime_acl_meter_index: .runtime_acl_meter_index, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        meter_metadata$meter_index <= runtime_acl_meter_index;
        acl_metadata$acl_copy <= runtime_acl_copy;
        fabric_metadata$reason_code <= runtime_acl_copy_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule acl_permit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged AclPermitRspT {pkt: pkt, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index, meter_metadata$meter_index: meter_metadata$meter_index, fabric_metadata$reason_code: fabric_metadata$reason_code, acl_metadata$acl_copy: acl_metadata$acl_copy};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== ACL_REDIRECT_ECMP ======

interface AclRedirectEcmp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkAclRedirectEcmp  (AclRedirectEcmp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) acl_metadata$acl_redirect <- mkReg(0);
  Reg#(Bit#(16)) acl_metadata$acl_nexthop <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_nexthop_type <- mkReg(0);
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(16)) meter_metadata$meter_index <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_copy <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule acl_redirect_ecmp_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged AclRedirectEcmpReqT {pkt: .pkt, runtime_acl_copy_reason: .runtime_acl_copy_reason, runtime_acl_meter_index: .runtime_acl_meter_index, runtime_acl_copy: .runtime_acl_copy, runtime_ecmp_index: .runtime_ecmp_index, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        acl_metadata$acl_redirect <= 'h1;
        acl_metadata$acl_nexthop <= runtime_ecmp_index;
        acl_metadata$acl_nexthop_type <= 'h1;
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        meter_metadata$meter_index <= runtime_acl_meter_index;
        acl_metadata$acl_copy <= runtime_acl_copy;
        fabric_metadata$reason_code <= runtime_acl_copy_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule acl_redirect_ecmp_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged AclRedirectEcmpRspT {pkt: pkt, meter_metadata$meter_index: meter_metadata$meter_index, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index, acl_metadata$acl_redirect: acl_metadata$acl_redirect, fabric_metadata$reason_code: fabric_metadata$reason_code, acl_metadata$acl_nexthop: acl_metadata$acl_nexthop, acl_metadata$acl_copy: acl_metadata$acl_copy, acl_metadata$acl_nexthop_type: acl_metadata$acl_nexthop_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== ACL_REDIRECT_NEXTHOP ======

interface AclRedirectNexthop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkAclRedirectNexthop  (AclRedirectNexthop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) acl_metadata$acl_redirect <- mkReg(0);
  Reg#(Bit#(16)) acl_metadata$acl_nexthop <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_nexthop_type <- mkReg(0);
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(16)) meter_metadata$meter_index <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_copy <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule acl_redirect_nexthop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged AclRedirectNexthopReqT {pkt: .pkt, runtime_acl_copy_reason: .runtime_acl_copy_reason, runtime_acl_meter_index: .runtime_acl_meter_index, runtime_acl_copy: .runtime_acl_copy, runtime_nexthop_index: .runtime_nexthop_index, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        acl_metadata$acl_redirect <= 'h1;
        acl_metadata$acl_nexthop <= runtime_nexthop_index;
        acl_metadata$acl_nexthop_type <= 'h0;
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        meter_metadata$meter_index <= runtime_acl_meter_index;
        acl_metadata$acl_copy <= runtime_acl_copy;
        fabric_metadata$reason_code <= runtime_acl_copy_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule acl_redirect_nexthop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged AclRedirectNexthopRspT {pkt: pkt, meter_metadata$meter_index: meter_metadata$meter_index, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index, acl_metadata$acl_redirect: acl_metadata$acl_redirect, fabric_metadata$reason_code: fabric_metadata$reason_code, acl_metadata$acl_nexthop: acl_metadata$acl_nexthop, acl_metadata$acl_copy: acl_metadata$acl_copy, acl_metadata$acl_nexthop_type: acl_metadata$acl_nexthop_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== ACL_STATS_UPDATE ======

interface AclStatsUpdate;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkAclStatsUpdate  (AclStatsUpdate);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule acl_stats_update_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged AclStatsUpdateReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule acl_stats_update_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged AclStatsUpdateRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== APPLY_COS_MARKING ======

interface ApplyCosMarking;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkApplyCosMarking  (ApplyCosMarking);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) qos_metadata$marked_cos <- mkReg(0);
  rule apply_cos_marking_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ApplyCosMarkingReqT {pkt: .pkt, runtime_cos: .runtime_cos}: begin
        qos_metadata$marked_cos <= runtime_cos;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule apply_cos_marking_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ApplyCosMarkingRspT {pkt: pkt, qos_metadata$marked_cos: qos_metadata$marked_cos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== APPLY_DSCP_MARKING ======

interface ApplyDscpMarking;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkApplyDscpMarking  (ApplyDscpMarking);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) qos_metadata$marked_dscp <- mkReg(0);
  rule apply_dscp_marking_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ApplyDscpMarkingReqT {pkt: .pkt, runtime_dscp: .runtime_dscp}: begin
        qos_metadata$marked_dscp <= runtime_dscp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule apply_dscp_marking_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ApplyDscpMarkingRspT {pkt: pkt, qos_metadata$marked_dscp: qos_metadata$marked_dscp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== APPLY_TC_MARKING ======

interface ApplyTcMarking;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkApplyTcMarking  (ApplyTcMarking);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) qos_metadata$marked_exp <- mkReg(0);
  rule apply_tc_marking_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ApplyTcMarkingReqT {pkt: .pkt, runtime_tc: .runtime_tc}: begin
        qos_metadata$marked_exp <= runtime_tc;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule apply_tc_marking_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ApplyTcMarkingRspT {pkt: pkt, qos_metadata$marked_exp: qos_metadata$marked_exp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== COMPUTE_LKP_IPV4_HASH ======

interface ComputeLkpIpv4Hash;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkComputeLkpIpv4Hash  (ComputeLkpIpv4Hash);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule compute_lkp_ipv4_hash_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ComputeLkpIpv4HashReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule compute_lkp_ipv4_hash_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ComputeLkpIpv4HashRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== COMPUTE_LKP_IPV6_HASH ======

interface ComputeLkpIpv6Hash;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkComputeLkpIpv6Hash  (ComputeLkpIpv6Hash);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule compute_lkp_ipv6_hash_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ComputeLkpIpv6HashReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule compute_lkp_ipv6_hash_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ComputeLkpIpv6HashRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== COMPUTE_LKP_NON_IP_HASH ======

interface ComputeLkpNonIpHash;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkComputeLkpNonIpHash  (ComputeLkpNonIpHash);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule compute_lkp_non_ip_hash_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ComputeLkpNonIpHashReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule compute_lkp_non_ip_hash_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ComputeLkpNonIpHashRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== COMPUTED_ONE_HASH ======

interface ComputedOneHash;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkComputedOneHash  (ComputedOneHash);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) hash_metadata$hash1 <- mkReg(0);
  Reg#(Bit#(13)) intrinsic_metadata$mcast_hash <- mkReg(0);
  Reg#(Bit#(16)) hash_metadata$entropy_hash <- mkReg(0);
  rule computed_one_hash_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ComputedOneHashReqT {pkt: .pkt, hash_metadata$hash2: .hash_metadata$hash2}: begin
        hash_metadata$hash1 <= hash_metadata$hash2;
        intrinsic_metadata$mcast_hash <= hash_metadata$hash2;
        hash_metadata$entropy_hash <= hash_metadata$hash2;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule computed_one_hash_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ComputedOneHashRspT {pkt: pkt, hash_metadata$entropy_hash: hash_metadata$entropy_hash, intrinsic_metadata$mcast_hash: intrinsic_metadata$mcast_hash, hash_metadata$hash1: hash_metadata$hash1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== COMPUTED_TWO_HASHES ======

interface ComputedTwoHashes;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkComputedTwoHashes  (ComputedTwoHashes);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(13)) intrinsic_metadata$mcast_hash <- mkReg(0);
  Reg#(Bit#(16)) hash_metadata$entropy_hash <- mkReg(0);
  rule computed_two_hashes_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ComputedTwoHashesReqT {pkt: .pkt, hash_metadata$hash1: .hash_metadata$hash1, hash_metadata$hash2: .hash_metadata$hash2}: begin
        intrinsic_metadata$mcast_hash <= hash_metadata$hash1;
        hash_metadata$entropy_hash <= hash_metadata$hash2;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule computed_two_hashes_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ComputedTwoHashesRspT {pkt: pkt, hash_metadata$entropy_hash: hash_metadata$entropy_hash, intrinsic_metadata$mcast_hash: intrinsic_metadata$mcast_hash};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== COPY_TO_CPU ======

interface CopyToCpu;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkCopyToCpu  (CopyToCpu);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule copy_to_cpu_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged CopyToCpuReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule copy_to_cpu_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged CopyToCpuRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== COPY_TO_CPU_WITH_REASON ======

interface CopyToCpuWithReason;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkCopyToCpuWithReason  (CopyToCpuWithReason);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule copy_to_cpu_with_reason_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged CopyToCpuWithReasonReqT {pkt: .pkt, runtime_reason_code: .runtime_reason_code}: begin
        fabric_metadata$reason_code <= runtime_reason_code;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule copy_to_cpu_with_reason_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged CopyToCpuWithReasonRspT {pkt: pkt, fabric_metadata$reason_code: fabric_metadata$reason_code};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== CPU_RX_REWRITE ======

interface CpuRxRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkCpuRxRewrite  (CpuRxRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) fabric_header$headerVersion <- mkReg(0);
  Reg#(Bit#(2)) fabric_header$packetVersion <- mkReg(0);
  Reg#(Bit#(1)) fabric_header$pad1 <- mkReg(0);
  Reg#(Bit#(3)) fabric_header$packetType <- mkReg(0);
  Reg#(Bit#(16)) fabric_header_cpu$ingressPort <- mkReg(0);
  Reg#(Bit#(16)) fabric_header_cpu$ingressIfindex <- mkReg(0);
  Reg#(Bit#(16)) fabric_header_cpu$ingressBd <- mkReg(0);
  Reg#(Bit#(16)) fabric_header_cpu$reasonCode <- mkReg(0);
  Reg#(Bit#(16)) fabric_payload_header$etherType <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule cpu_rx_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged CpuRxRewriteReqT {pkt: .pkt, ingress_metadata$bd: .ingress_metadata$bd, fabric_metadata$reason_code: .fabric_metadata$reason_code, ingress_metadata$ingress_port: .ingress_metadata$ingress_port, ingress_metadata$ifindex: .ingress_metadata$ifindex, ethernet$etherType: .ethernet$etherType}: begin
        fabric_header$headerVersion <= 'h0;
        fabric_header$packetVersion <= 'h0;
        fabric_header$pad1 <= 'h0;
        fabric_header$packetType <= 'h5;
        fabric_header_cpu$ingressPort <= ingress_metadata$ingress_port;
        fabric_header_cpu$ingressIfindex <= ingress_metadata$ifindex;
        fabric_header_cpu$ingressBd <= ingress_metadata$bd;
        fabric_header_cpu$reasonCode <= fabric_metadata$reason_code;
        fabric_payload_header$etherType <= ethernet$etherType;
        ethernet$etherType <= 'h9000;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule cpu_rx_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged CpuRxRewriteRspT {pkt: pkt, fabric_header$packetType: fabric_header$packetType, fabric_header_cpu$reasonCode: fabric_header_cpu$reasonCode, fabric_header_cpu$ingressPort: fabric_header_cpu$ingressPort, fabric_header_cpu$ingressIfindex: fabric_header_cpu$ingressIfindex, fabric_payload_header$etherType: fabric_payload_header$etherType, fabric_header_cpu$ingressBd: fabric_header_cpu$ingressBd, fabric_header$headerVersion: fabric_header$headerVersion, fabric_header$packetVersion: fabric_header$packetVersion, ethernet$etherType: ethernet$etherType, fabric_header$pad1: fabric_header$pad1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_GENV_INNER_IPV4 ======

interface DecapGenvInnerIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapGenvInnerIpv4  (DecapGenvInnerIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_genv_inner_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapGenvInnerIpv4ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_genv_inner_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapGenvInnerIpv4RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_GENV_INNER_IPV6 ======

interface DecapGenvInnerIpv6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapGenvInnerIpv6  (DecapGenvInnerIpv6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_genv_inner_ipv6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapGenvInnerIpv6ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_genv_inner_ipv6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapGenvInnerIpv6RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_GENV_INNER_NON_IP ======

interface DecapGenvInnerNonIp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapGenvInnerNonIp  (DecapGenvInnerNonIp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_genv_inner_non_ip_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapGenvInnerNonIpReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_genv_inner_non_ip_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapGenvInnerNonIpRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_GRE_INNER_IPV4 ======

interface DecapGreInnerIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapGreInnerIpv4  (DecapGreInnerIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_gre_inner_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapGreInnerIpv4ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_gre_inner_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapGreInnerIpv4RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_GRE_INNER_IPV6 ======

interface DecapGreInnerIpv6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapGreInnerIpv6  (DecapGreInnerIpv6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_gre_inner_ipv6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapGreInnerIpv6ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_gre_inner_ipv6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapGreInnerIpv6RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_GRE_INNER_NON_IP ======

interface DecapGreInnerNonIp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapGreInnerNonIp  (DecapGreInnerNonIp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_gre_inner_non_ip_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapGreInnerNonIpReqT {pkt: .pkt, gre$proto: .gre$proto}: begin
        ethernet$etherType <= gre$proto;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_gre_inner_non_ip_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapGreInnerNonIpRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_INNER_ICMP ======

interface DecapInnerIcmp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapInnerIcmp  (DecapInnerIcmp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_inner_icmp_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapInnerIcmpReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_inner_icmp_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapInnerIcmpRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_INNER_TCP ======

interface DecapInnerTcp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapInnerTcp  (DecapInnerTcp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_inner_tcp_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapInnerTcpReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_inner_tcp_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapInnerTcpRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_INNER_UDP ======

interface DecapInnerUdp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapInnerUdp  (DecapInnerUdp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_inner_udp_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapInnerUdpReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_inner_udp_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapInnerUdpRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_INNER_UNKNOWN ======

interface DecapInnerUnknown;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapInnerUnknown  (DecapInnerUnknown);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_inner_unknown_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapInnerUnknownReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_inner_unknown_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapInnerUnknownRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_IP_INNER_IPV4 ======

interface DecapIpInnerIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapIpInnerIpv4  (DecapIpInnerIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_ip_inner_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapIpInnerIpv4ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_ip_inner_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapIpInnerIpv4RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_IP_INNER_IPV6 ======

interface DecapIpInnerIpv6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapIpInnerIpv6  (DecapIpInnerIpv6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_ip_inner_ipv6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapIpInnerIpv6ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_ip_inner_ipv6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapIpInnerIpv6RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_IPV4_POP1 ======

interface DecapMplsInnerEthernetIpv4Pop1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetIpv4Pop1  (DecapMplsInnerEthernetIpv4Pop1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_ipv4_pop1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetIpv4Pop1ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_ipv4_pop1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetIpv4Pop1RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_IPV4_POP2 ======

interface DecapMplsInnerEthernetIpv4Pop2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetIpv4Pop2  (DecapMplsInnerEthernetIpv4Pop2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_ipv4_pop2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetIpv4Pop2ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_ipv4_pop2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetIpv4Pop2RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_IPV4_POP3 ======

interface DecapMplsInnerEthernetIpv4Pop3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetIpv4Pop3  (DecapMplsInnerEthernetIpv4Pop3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_ipv4_pop3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetIpv4Pop3ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_ipv4_pop3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetIpv4Pop3RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_IPV6_POP1 ======

interface DecapMplsInnerEthernetIpv6Pop1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetIpv6Pop1  (DecapMplsInnerEthernetIpv6Pop1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_ipv6_pop1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetIpv6Pop1ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_ipv6_pop1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetIpv6Pop1RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_IPV6_POP2 ======

interface DecapMplsInnerEthernetIpv6Pop2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetIpv6Pop2  (DecapMplsInnerEthernetIpv6Pop2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_ipv6_pop2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetIpv6Pop2ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_ipv6_pop2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetIpv6Pop2RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_IPV6_POP3 ======

interface DecapMplsInnerEthernetIpv6Pop3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetIpv6Pop3  (DecapMplsInnerEthernetIpv6Pop3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_ipv6_pop3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetIpv6Pop3ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_ipv6_pop3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetIpv6Pop3RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_NON_IP_POP1 ======

interface DecapMplsInnerEthernetNonIpPop1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetNonIpPop1  (DecapMplsInnerEthernetNonIpPop1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_non_ip_pop1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetNonIpPop1ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_non_ip_pop1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetNonIpPop1RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_NON_IP_POP2 ======

interface DecapMplsInnerEthernetNonIpPop2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetNonIpPop2  (DecapMplsInnerEthernetNonIpPop2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_non_ip_pop2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetNonIpPop2ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_non_ip_pop2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetNonIpPop2RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_ETHERNET_NON_IP_POP3 ======

interface DecapMplsInnerEthernetNonIpPop3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerEthernetNonIpPop3  (DecapMplsInnerEthernetNonIpPop3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_mpls_inner_ethernet_non_ip_pop3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerEthernetNonIpPop3ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ethernet_non_ip_pop3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerEthernetNonIpPop3RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_IPV4_POP1 ======

interface DecapMplsInnerIpv4Pop1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerIpv4Pop1  (DecapMplsInnerIpv4Pop1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_mpls_inner_ipv4_pop1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerIpv4Pop1ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ipv4_pop1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerIpv4Pop1RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_IPV4_POP2 ======

interface DecapMplsInnerIpv4Pop2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerIpv4Pop2  (DecapMplsInnerIpv4Pop2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_mpls_inner_ipv4_pop2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerIpv4Pop2ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ipv4_pop2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerIpv4Pop2RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_IPV4_POP3 ======

interface DecapMplsInnerIpv4Pop3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerIpv4Pop3  (DecapMplsInnerIpv4Pop3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_mpls_inner_ipv4_pop3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerIpv4Pop3ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ipv4_pop3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerIpv4Pop3RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_IPV6_POP1 ======

interface DecapMplsInnerIpv6Pop1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerIpv6Pop1  (DecapMplsInnerIpv6Pop1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_mpls_inner_ipv6_pop1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerIpv6Pop1ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ipv6_pop1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerIpv6Pop1RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_IPV6_POP2 ======

interface DecapMplsInnerIpv6Pop2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerIpv6Pop2  (DecapMplsInnerIpv6Pop2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_mpls_inner_ipv6_pop2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerIpv6Pop2ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ipv6_pop2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerIpv6Pop2RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_MPLS_INNER_IPV6_POP3 ======

interface DecapMplsInnerIpv6Pop3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapMplsInnerIpv6Pop3  (DecapMplsInnerIpv6Pop3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule decap_mpls_inner_ipv6_pop3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapMplsInnerIpv6Pop3ReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_mpls_inner_ipv6_pop3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapMplsInnerIpv6Pop3RspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_NVGRE_INNER_IPV4 ======

interface DecapNvgreInnerIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapNvgreInnerIpv4  (DecapNvgreInnerIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_nvgre_inner_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapNvgreInnerIpv4ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_nvgre_inner_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapNvgreInnerIpv4RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_NVGRE_INNER_IPV6 ======

interface DecapNvgreInnerIpv6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapNvgreInnerIpv6  (DecapNvgreInnerIpv6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_nvgre_inner_ipv6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapNvgreInnerIpv6ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_nvgre_inner_ipv6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapNvgreInnerIpv6RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_NVGRE_INNER_NON_IP ======

interface DecapNvgreInnerNonIp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapNvgreInnerNonIp  (DecapNvgreInnerNonIp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_nvgre_inner_non_ip_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapNvgreInnerNonIpReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_nvgre_inner_non_ip_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapNvgreInnerNonIpRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_VXLAN_INNER_IPV4 ======

interface DecapVxlanInnerIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapVxlanInnerIpv4  (DecapVxlanInnerIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_vxlan_inner_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapVxlanInnerIpv4ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_vxlan_inner_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapVxlanInnerIpv4RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_VXLAN_INNER_IPV6 ======

interface DecapVxlanInnerIpv6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapVxlanInnerIpv6  (DecapVxlanInnerIpv6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_vxlan_inner_ipv6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapVxlanInnerIpv6ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_vxlan_inner_ipv6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapVxlanInnerIpv6RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DECAP_VXLAN_INNER_NON_IP ======

interface DecapVxlanInnerNonIp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDecapVxlanInnerNonIp  (DecapVxlanInnerNonIp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule decap_vxlan_inner_non_ip_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DecapVxlanInnerNonIpReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule decap_vxlan_inner_non_ip_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DecapVxlanInnerNonIpRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DMAC_DROP ======

interface DmacDrop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDmacDrop  (DmacDrop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule dmac_drop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DmacDropReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule dmac_drop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DmacDropRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DMAC_HIT ======

interface DmacHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDmacHit  (DmacHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  rule dmac_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DmacHitReqT {pkt: .pkt, runtime_ifindex: .runtime_ifindex}: begin
        ingress_metadata$egress_ifindex <= runtime_ifindex;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule dmac_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DmacHitRspT {pkt: pkt, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DMAC_MISS ======

interface DmacMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDmacMiss  (DmacMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule dmac_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DmacMissReqT {pkt: .pkt}: begin
        ingress_metadata$egress_ifindex <= 'hffff;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule dmac_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DmacMissRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DMAC_MULTICAST_HIT ======

interface DmacMulticastHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDmacMulticastHit  (DmacMulticastHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule dmac_multicast_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DmacMulticastHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index}: begin
        intrinsic_metadata$mcast_grp <= runtime_mc_index;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule dmac_multicast_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DmacMulticastHitRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DMAC_REDIRECT_ECMP ======

interface DmacRedirectEcmp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDmacRedirectEcmp  (DmacRedirectEcmp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l2_metadata$l2_redirect <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$l2_nexthop <- mkReg(0);
  Reg#(Bit#(1)) l2_metadata$l2_nexthop_type <- mkReg(0);
  rule dmac_redirect_ecmp_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DmacRedirectEcmpReqT {pkt: .pkt, runtime_ecmp_index: .runtime_ecmp_index}: begin
        l2_metadata$l2_redirect <= 'h1;
        l2_metadata$l2_nexthop <= runtime_ecmp_index;
        l2_metadata$l2_nexthop_type <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule dmac_redirect_ecmp_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DmacRedirectEcmpRspT {pkt: pkt, l2_metadata$l2_redirect: l2_metadata$l2_redirect, l2_metadata$l2_nexthop: l2_metadata$l2_nexthop, l2_metadata$l2_nexthop_type: l2_metadata$l2_nexthop_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DMAC_REDIRECT_NEXTHOP ======

interface DmacRedirectNexthop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDmacRedirectNexthop  (DmacRedirectNexthop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l2_metadata$l2_redirect <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$l2_nexthop <- mkReg(0);
  Reg#(Bit#(1)) l2_metadata$l2_nexthop_type <- mkReg(0);
  rule dmac_redirect_nexthop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DmacRedirectNexthopReqT {pkt: .pkt, runtime_nexthop_index: .runtime_nexthop_index}: begin
        l2_metadata$l2_redirect <= 'h1;
        l2_metadata$l2_nexthop <= runtime_nexthop_index;
        l2_metadata$l2_nexthop_type <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule dmac_redirect_nexthop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DmacRedirectNexthopRspT {pkt: pkt, l2_metadata$l2_redirect: l2_metadata$l2_redirect, l2_metadata$l2_nexthop: l2_metadata$l2_nexthop, l2_metadata$l2_nexthop_type: l2_metadata$l2_nexthop_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DROP_PACKET ======

interface DropPacket;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDropPacket  (DropPacket);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule drop_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DropPacketReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule drop_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DropPacketRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DROP_PACKET_WITH_REASON ======

interface DropPacketWithReason;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDropPacketWithReason  (DropPacketWithReason);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule drop_packet_with_reason_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DropPacketWithReasonReqT {pkt: .pkt, runtime_drop_reason: .runtime_drop_reason}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule drop_packet_with_reason_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DropPacketWithReasonRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== DROP_STATS_UPDATE ======

interface DropStatsUpdate;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkDropStatsUpdate  (DropStatsUpdate);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule drop_stats_update_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged DropStatsUpdateReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule drop_stats_update_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged DropStatsUpdateRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== EGRESS_FILTER_CHECK ======

interface EgressFilterCheck;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkEgressFilterCheck  (EgressFilterCheck);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule egress_filter_check_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged EgressFilterCheckReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule egress_filter_check_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged EgressFilterCheckRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== EGRESS_MIRROR ======

interface EgressMirror;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkEgressMirror  (EgressMirror);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) i2e_metadata$mirror_session_id <- mkReg(0);
  rule egress_mirror_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged EgressMirrorReqT {pkt: .pkt, runtime_session_id: .runtime_session_id}: begin
        i2e_metadata$mirror_session_id <= runtime_session_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule egress_mirror_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged EgressMirrorRspT {pkt: pkt, i2e_metadata$mirror_session_id: i2e_metadata$mirror_session_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== EGRESS_MIRROR_DROP ======

interface EgressMirrorDrop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkEgressMirrorDrop  (EgressMirrorDrop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) i2e_metadata$mirror_session_id <- mkReg(0);
  rule egress_mirror_drop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged EgressMirrorDropReqT {pkt: .pkt, runtime_session_id: .runtime_session_id}: begin
        i2e_metadata$mirror_session_id <= runtime_session_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule egress_mirror_drop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged EgressMirrorDropRspT {pkt: pkt, i2e_metadata$mirror_session_id: i2e_metadata$mirror_session_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== EGRESS_PORT_TYPE_CPU ======

interface EgressPortTypeCpu;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkEgressPortTypeCpu  (EgressPortTypeCpu);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) egress_metadata$port_type <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$ifindex <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  rule egress_port_type_cpu_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged EgressPortTypeCpuReqT {pkt: .pkt, runtime_ifindex: .runtime_ifindex}: begin
        egress_metadata$port_type <= 'h2;
        egress_metadata$ifindex <= runtime_ifindex;
        tunnel_metadata$egress_tunnel_type <= 'h10;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule egress_port_type_cpu_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged EgressPortTypeCpuRspT {pkt: pkt, egress_metadata$ifindex: egress_metadata$ifindex, egress_metadata$port_type: egress_metadata$port_type, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== EGRESS_PORT_TYPE_FABRIC ======

interface EgressPortTypeFabric;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkEgressPortTypeFabric  (EgressPortTypeFabric);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) egress_metadata$port_type <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$ifindex <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  rule egress_port_type_fabric_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged EgressPortTypeFabricReqT {pkt: .pkt, runtime_ifindex: .runtime_ifindex}: begin
        egress_metadata$port_type <= 'h1;
        egress_metadata$ifindex <= runtime_ifindex;
        tunnel_metadata$egress_tunnel_type <= 'hf;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule egress_port_type_fabric_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged EgressPortTypeFabricRspT {pkt: pkt, egress_metadata$ifindex: egress_metadata$ifindex, egress_metadata$port_type: egress_metadata$port_type, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== EGRESS_PORT_TYPE_NORMAL ======

interface EgressPortTypeNormal;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkEgressPortTypeNormal  (EgressPortTypeNormal);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) egress_metadata$port_type <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$ifindex <- mkReg(0);
  rule egress_port_type_normal_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged EgressPortTypeNormalReqT {pkt: .pkt, runtime_ifindex: .runtime_ifindex}: begin
        egress_metadata$port_type <= 'h0;
        egress_metadata$ifindex <= runtime_ifindex;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule egress_port_type_normal_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged EgressPortTypeNormalRspT {pkt: pkt, egress_metadata$ifindex: egress_metadata$ifindex, egress_metadata$port_type: egress_metadata$port_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== EGRESS_REDIRECT_TO_CPU ======

interface EgressRedirectToCpu;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkEgressRedirectToCpu  (EgressRedirectToCpu);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule egress_redirect_to_cpu_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged EgressRedirectToCpuReqT {pkt: .pkt, runtime_reason_code: .runtime_reason_code}: begin
        fabric_metadata$reason_code <= runtime_reason_code;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule egress_redirect_to_cpu_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged EgressRedirectToCpuRspT {pkt: pkt, fabric_metadata$reason_code: fabric_metadata$reason_code};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== FABRIC_MULTICAST_REWRITE ======

interface FabricMulticastRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkFabricMulticastRewrite  (FabricMulticastRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) fabric_header$headerVersion <- mkReg(0);
  Reg#(Bit#(2)) fabric_header$packetVersion <- mkReg(0);
  Reg#(Bit#(1)) fabric_header$pad1 <- mkReg(0);
  Reg#(Bit#(3)) fabric_header$packetType <- mkReg(0);
  Reg#(Bit#(8)) fabric_header$dstDevice <- mkReg(0);
  Reg#(Bit#(16)) fabric_header$dstPortOrGroup <- mkReg(0);
  Reg#(Bit#(16)) fabric_header_multicast$ingressIfindex <- mkReg(0);
  Reg#(Bit#(16)) fabric_header_multicast$ingressBd <- mkReg(0);
  Reg#(Bit#(1)) fabric_header_multicast$tunnelTerminate <- mkReg(0);
  Reg#(Bit#(1)) fabric_header_multicast$routed <- mkReg(0);
  Reg#(Bit#(1)) fabric_header_multicast$outerRouted <- mkReg(0);
  Reg#(Bit#(5)) fabric_header_multicast$ingressTunnelType <- mkReg(0);
  Reg#(Bit#(16)) fabric_header_multicast$mcastGrp <- mkReg(0);
  Reg#(Bit#(16)) fabric_payload_header$etherType <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule fabric_multicast_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged FabricMulticastRewriteReqT {pkt: .pkt, multicast_metadata$mcast_grp: .multicast_metadata$mcast_grp, ingress_metadata$bd: .ingress_metadata$bd, tunnel_metadata$ingress_tunnel_type: .tunnel_metadata$ingress_tunnel_type, l3_metadata$routed: .l3_metadata$routed, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, ingress_metadata$ifindex: .ingress_metadata$ifindex, ethernet$etherType: .ethernet$etherType, l3_metadata$outer_routed: .l3_metadata$outer_routed, runtime_fabric_mgid: .runtime_fabric_mgid}: begin
        fabric_header$headerVersion <= 'h0;
        fabric_header$packetVersion <= 'h0;
        fabric_header$pad1 <= 'h0;
        fabric_header$packetType <= 'h2;
        fabric_header$dstDevice <= 'h7f;
        fabric_header$dstPortOrGroup <= runtime_fabric_mgid;
        fabric_header_multicast$ingressIfindex <= ingress_metadata$ifindex;
        fabric_header_multicast$ingressBd <= ingress_metadata$bd;
        fabric_header_multicast$tunnelTerminate <= tunnel_metadata$tunnel_terminate;
        fabric_header_multicast$routed <= l3_metadata$routed;
        fabric_header_multicast$outerRouted <= l3_metadata$outer_routed;
        fabric_header_multicast$ingressTunnelType <= tunnel_metadata$ingress_tunnel_type;
        fabric_header_multicast$mcastGrp <= multicast_metadata$mcast_grp;
        fabric_payload_header$etherType <= ethernet$etherType;
        ethernet$etherType <= 'h9000;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule fabric_multicast_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged FabricMulticastRewriteRspT {pkt: pkt, fabric_header$packetType: fabric_header$packetType, fabric_header_multicast$tunnelTerminate: fabric_header_multicast$tunnelTerminate, fabric_header_multicast$routed: fabric_header_multicast$routed, fabric_header_multicast$ingressTunnelType: fabric_header_multicast$ingressTunnelType, fabric_header$dstDevice: fabric_header$dstDevice, fabric_header_multicast$outerRouted: fabric_header_multicast$outerRouted, fabric_header_multicast$ingressIfindex: fabric_header_multicast$ingressIfindex, fabric_header$dstPortOrGroup: fabric_header$dstPortOrGroup, fabric_payload_header$etherType: fabric_payload_header$etherType, fabric_header_multicast$ingressBd: fabric_header_multicast$ingressBd, fabric_header_multicast$mcastGrp: fabric_header_multicast$mcastGrp, fabric_header$pad1: fabric_header$pad1, fabric_header$packetVersion: fabric_header$packetVersion, ethernet$etherType: ethernet$etherType, fabric_header$headerVersion: fabric_header$headerVersion};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== FABRIC_REWRITE ======

interface FabricRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkFabricRewrite  (FabricRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  rule fabric_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged FabricRewriteReqT {pkt: .pkt, runtime_tunnel_index: .runtime_tunnel_index}: begin
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule fabric_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged FabricRewriteRspT {pkt: pkt, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== FABRIC_UNICAST_REWRITE ======

interface FabricUnicastRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkFabricUnicastRewrite  (FabricUnicastRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) fabric_header$headerVersion <- mkReg(0);
  Reg#(Bit#(2)) fabric_header$packetVersion <- mkReg(0);
  Reg#(Bit#(1)) fabric_header$pad1 <- mkReg(0);
  Reg#(Bit#(3)) fabric_header$packetType <- mkReg(0);
  Reg#(Bit#(8)) fabric_header$dstDevice <- mkReg(0);
  Reg#(Bit#(16)) fabric_header$dstPortOrGroup <- mkReg(0);
  Reg#(Bit#(1)) fabric_header_unicast$tunnelTerminate <- mkReg(0);
  Reg#(Bit#(1)) fabric_header_unicast$routed <- mkReg(0);
  Reg#(Bit#(1)) fabric_header_unicast$outerRouted <- mkReg(0);
  Reg#(Bit#(5)) fabric_header_unicast$ingressTunnelType <- mkReg(0);
  Reg#(Bit#(16)) fabric_header_unicast$nexthopIndex <- mkReg(0);
  Reg#(Bit#(16)) fabric_payload_header$etherType <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule fabric_unicast_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged FabricUnicastRewriteReqT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, tunnel_metadata$ingress_tunnel_type: .tunnel_metadata$ingress_tunnel_type, l3_metadata$routed: .l3_metadata$routed, fabric_metadata$dst_device: .fabric_metadata$dst_device, fabric_metadata$dst_port: .fabric_metadata$dst_port, ethernet$etherType: .ethernet$etherType, l3_metadata$outer_routed: .l3_metadata$outer_routed}: begin
        fabric_header$headerVersion <= 'h0;
        fabric_header$packetVersion <= 'h0;
        fabric_header$pad1 <= 'h0;
        fabric_header$packetType <= 'h1;
        fabric_header$dstDevice <= fabric_metadata$dst_device;
        fabric_header$dstPortOrGroup <= fabric_metadata$dst_port;
        fabric_header_unicast$tunnelTerminate <= tunnel_metadata$tunnel_terminate;
        fabric_header_unicast$routed <= l3_metadata$routed;
        fabric_header_unicast$outerRouted <= l3_metadata$outer_routed;
        fabric_header_unicast$ingressTunnelType <= tunnel_metadata$ingress_tunnel_type;
        fabric_header_unicast$nexthopIndex <= l3_metadata$nexthop_index;
        fabric_payload_header$etherType <= ethernet$etherType;
        ethernet$etherType <= 'h9000;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule fabric_unicast_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged FabricUnicastRewriteRspT {pkt: pkt, fabric_header$packetType: fabric_header$packetType, fabric_header_unicast$outerRouted: fabric_header_unicast$outerRouted, fabric_header_unicast$tunnelTerminate: fabric_header_unicast$tunnelTerminate, fabric_payload_header$etherType: fabric_payload_header$etherType, fabric_header$dstDevice: fabric_header$dstDevice, fabric_header_unicast$ingressTunnelType: fabric_header_unicast$ingressTunnelType, fabric_header$dstPortOrGroup: fabric_header$dstPortOrGroup, fabric_header_unicast$nexthopIndex: fabric_header_unicast$nexthopIndex, fabric_header_unicast$routed: fabric_header_unicast$routed, fabric_header$pad1: fabric_header$pad1, fabric_header$packetVersion: fabric_header$packetVersion, ethernet$etherType: ethernet$etherType, fabric_header$headerVersion: fabric_header$headerVersion};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== FIB_HIT_ECMP ======

interface FibHitEcmp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkFibHitEcmp  (FibHitEcmp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$fib_hit <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$fib_nexthop <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$fib_nexthop_type <- mkReg(0);
  rule fib_hit_ecmp_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged FibHitEcmpReqT {pkt: .pkt, runtime_ecmp_index: .runtime_ecmp_index}: begin
        l3_metadata$fib_hit <= 'h1;
        l3_metadata$fib_nexthop <= runtime_ecmp_index;
        l3_metadata$fib_nexthop_type <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule fib_hit_ecmp_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged FibHitEcmpRspT {pkt: pkt, l3_metadata$fib_nexthop: l3_metadata$fib_nexthop, l3_metadata$fib_hit: l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: l3_metadata$fib_nexthop_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== FIB_HIT_NEXTHOP ======

interface FibHitNexthop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkFibHitNexthop  (FibHitNexthop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$fib_hit <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$fib_nexthop <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$fib_nexthop_type <- mkReg(0);
  rule fib_hit_nexthop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged FibHitNexthopReqT {pkt: .pkt, runtime_nexthop_index: .runtime_nexthop_index}: begin
        l3_metadata$fib_hit <= 'h1;
        l3_metadata$fib_nexthop <= runtime_nexthop_index;
        l3_metadata$fib_nexthop_type <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule fib_hit_nexthop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged FibHitNexthopRspT {pkt: pkt, l3_metadata$fib_nexthop: l3_metadata$fib_nexthop, l3_metadata$fib_hit: l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: l3_metadata$fib_nexthop_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== FORWARD_MPLS ======

interface ForwardMpls;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkForwardMpls  (ForwardMpls);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) l3_metadata$fib_nexthop <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$fib_nexthop_type <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$fib_hit <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  rule forward_mpls_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged ForwardMplsReqT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, runtime_nexthop_index: .runtime_nexthop_index}: begin
        l3_metadata$fib_nexthop <= runtime_nexthop_index;
        l3_metadata$fib_nexthop_type <= 'h0;
        l3_metadata$fib_hit <= 'h1;
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule forward_mpls_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged ForwardMplsRspT {pkt: pkt, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l3_metadata$fib_nexthop: l3_metadata$fib_nexthop, l3_metadata$fib_hit: l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: l3_metadata$fib_nexthop_type, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== GENERATE_LEARN_NOTIFY ======

interface GenerateLearnNotify;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkGenerateLearnNotify  (GenerateLearnNotify);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule generate_learn_notify_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged GenerateLearnNotifyReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule generate_learn_notify_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged GenerateLearnNotifyRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_IPV4_ICMP_REWRITE ======

interface InnerIpv4IcmpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerIpv4IcmpRewrite  (InnerIpv4IcmpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) egress_metadata$payload_length <- mkReg(0);
  Reg#(Bit#(8)) tunnel_metadata$inner_ip_proto <- mkReg(0);
  rule inner_ipv4_icmp_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerIpv4IcmpRewriteReqT {pkt: .pkt, ipv4$totalLen: .ipv4$totalLen}: begin
        egress_metadata$payload_length <= ipv4$totalLen;
        tunnel_metadata$inner_ip_proto <= 'h4;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_ipv4_icmp_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerIpv4IcmpRewriteRspT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: egress_metadata$payload_length};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_IPV4_TCP_REWRITE ======

interface InnerIpv4TcpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerIpv4TcpRewrite  (InnerIpv4TcpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) egress_metadata$payload_length <- mkReg(0);
  Reg#(Bit#(8)) tunnel_metadata$inner_ip_proto <- mkReg(0);
  rule inner_ipv4_tcp_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerIpv4TcpRewriteReqT {pkt: .pkt, ipv4$totalLen: .ipv4$totalLen}: begin
        egress_metadata$payload_length <= ipv4$totalLen;
        tunnel_metadata$inner_ip_proto <= 'h4;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_ipv4_tcp_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerIpv4TcpRewriteRspT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: egress_metadata$payload_length};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_IPV4_UDP_REWRITE ======

interface InnerIpv4UdpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerIpv4UdpRewrite  (InnerIpv4UdpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) egress_metadata$payload_length <- mkReg(0);
  Reg#(Bit#(8)) tunnel_metadata$inner_ip_proto <- mkReg(0);
  rule inner_ipv4_udp_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerIpv4UdpRewriteReqT {pkt: .pkt, ipv4$totalLen: .ipv4$totalLen}: begin
        egress_metadata$payload_length <= ipv4$totalLen;
        tunnel_metadata$inner_ip_proto <= 'h4;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_ipv4_udp_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerIpv4UdpRewriteRspT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: egress_metadata$payload_length};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_IPV4_UNKNOWN_REWRITE ======

interface InnerIpv4UnknownRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerIpv4UnknownRewrite  (InnerIpv4UnknownRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) egress_metadata$payload_length <- mkReg(0);
  Reg#(Bit#(8)) tunnel_metadata$inner_ip_proto <- mkReg(0);
  rule inner_ipv4_unknown_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerIpv4UnknownRewriteReqT {pkt: .pkt, ipv4$totalLen: .ipv4$totalLen}: begin
        egress_metadata$payload_length <= ipv4$totalLen;
        tunnel_metadata$inner_ip_proto <= 'h4;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_ipv4_unknown_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerIpv4UnknownRewriteRspT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: egress_metadata$payload_length};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_IPV6_ICMP_REWRITE ======

interface InnerIpv6IcmpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerIpv6IcmpRewrite  (InnerIpv6IcmpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) tunnel_metadata$inner_ip_proto <- mkReg(0);
  rule inner_ipv6_icmp_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerIpv6IcmpRewriteReqT {pkt: .pkt}: begin
        tunnel_metadata$inner_ip_proto <= 'h29;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_ipv6_icmp_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerIpv6IcmpRewriteRspT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_IPV6_TCP_REWRITE ======

interface InnerIpv6TcpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerIpv6TcpRewrite  (InnerIpv6TcpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) tunnel_metadata$inner_ip_proto <- mkReg(0);
  rule inner_ipv6_tcp_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerIpv6TcpRewriteReqT {pkt: .pkt}: begin
        tunnel_metadata$inner_ip_proto <= 'h29;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_ipv6_tcp_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerIpv6TcpRewriteRspT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_IPV6_UDP_REWRITE ======

interface InnerIpv6UdpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerIpv6UdpRewrite  (InnerIpv6UdpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) tunnel_metadata$inner_ip_proto <- mkReg(0);
  rule inner_ipv6_udp_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerIpv6UdpRewriteReqT {pkt: .pkt}: begin
        tunnel_metadata$inner_ip_proto <= 'h29;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_ipv6_udp_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerIpv6UdpRewriteRspT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_IPV6_UNKNOWN_REWRITE ======

interface InnerIpv6UnknownRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerIpv6UnknownRewrite  (InnerIpv6UnknownRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) tunnel_metadata$inner_ip_proto <- mkReg(0);
  rule inner_ipv6_unknown_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerIpv6UnknownRewriteReqT {pkt: .pkt}: begin
        tunnel_metadata$inner_ip_proto <= 'h29;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_ipv6_unknown_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerIpv6UnknownRewriteRspT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_NON_IP_REWRITE ======

interface InnerNonIpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerNonIpRewrite  (InnerNonIpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule inner_non_ip_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerNonIpRewriteReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_non_ip_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerNonIpRewriteRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INNER_REPLICA_FROM_RID ======

interface InnerReplicaFromRid;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkInnerReplicaFromRid  (InnerReplicaFromRid);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$replica <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$inner_replica <- mkReg(0);
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  Reg#(Bit#(4)) tunnel_metadata$egress_header_count <- mkReg(0);
  rule inner_replica_from_rid_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged InnerReplicaFromRidReqT {pkt: .pkt, l3_metadata$routed: .l3_metadata$routed, runtime_tunnel_index: .runtime_tunnel_index, runtime_tunnel_type: .runtime_tunnel_type, runtime_bd: .runtime_bd, runtime_header_count: .runtime_header_count}: begin
        egress_metadata$bd <= runtime_bd;
        multicast_metadata$replica <= 'h1;
        multicast_metadata$inner_replica <= 'h1;
        egress_metadata$routed <= l3_metadata$routed;
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        tunnel_metadata$egress_tunnel_type <= runtime_tunnel_type;
        tunnel_metadata$egress_header_count <= runtime_header_count;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule inner_replica_from_rid_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged InnerReplicaFromRidRspT {pkt: pkt, multicast_metadata$replica: multicast_metadata$replica, multicast_metadata$inner_replica: multicast_metadata$inner_replica, tunnel_metadata$egress_header_count: tunnel_metadata$egress_header_count, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type, egress_metadata$bd: egress_metadata$bd, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index, egress_metadata$routed: egress_metadata$routed};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_ADD_UPDATE_VXLAN_GPE_IPV4 ======

interface IntAddUpdateVxlanGpeIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntAddUpdateVxlanGpeIpv4  (IntAddUpdateVxlanGpeIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) vxlan_gpe_int_header$int_type <- mkReg(0);
  Reg#(Bit#(8)) vxlan_gpe_int_header$next_proto <- mkReg(0);
  Reg#(Bit#(8)) vxlan_gpe$next_proto <- mkReg(0);
  Reg#(Bit#(8)) vxlan_gpe_int_header$len <- mkReg(0);
  rule int_add_update_vxlan_gpe_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntAddUpdateVxlanGpeIpv4ReqT {pkt: .pkt, int_metadata$gpe_int_hdr_len8: .int_metadata$gpe_int_hdr_len8, int_metadata$insert_byte_cnt: .int_metadata$insert_byte_cnt}: begin
        vxlan_gpe_int_header$int_type <= 'h1;
        vxlan_gpe_int_header$next_proto <= 'h3;
        vxlan_gpe$next_proto <= 'h5;
        vxlan_gpe_int_header$len <= int_metadata$gpe_int_hdr_len8;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_add_update_vxlan_gpe_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntAddUpdateVxlanGpeIpv4RspT {pkt: pkt, vxlan_gpe$next_proto: vxlan_gpe$next_proto, vxlan_gpe_int_header$len: vxlan_gpe_int_header$len, vxlan_gpe_int_header$next_proto: vxlan_gpe_int_header$next_proto, vxlan_gpe_int_header$int_type: vxlan_gpe_int_header$int_type, udp$length_: udp$length_, ipv4$totalLen: ipv4$totalLen};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_NO_SINK ======

interface IntNoSink;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntNoSink  (IntNoSink);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_metadata_i2e$sink <- mkReg(0);
  rule int_no_sink_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntNoSinkReqT {pkt: .pkt}: begin
        int_metadata_i2e$sink <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_no_sink_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntNoSinkRspT {pkt: pkt, int_metadata_i2e$sink: int_metadata_i2e$sink};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_RESET ======

interface IntReset;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntReset  (IntReset);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(32)) int_metadata$switch_id <- mkReg(0);
  Reg#(Bit#(16)) int_metadata$insert_byte_cnt <- mkReg(0);
  Reg#(Bit#(8)) int_metadata$insert_cnt <- mkReg(0);
  Reg#(Bit#(8)) int_metadata$gpe_int_hdr_len8 <- mkReg(0);
  Reg#(Bit#(16)) int_metadata$gpe_int_hdr_len <- mkReg(0);
  Reg#(Bit#(16)) int_metadata$instruction_cnt <- mkReg(0);
  rule int_reset_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntResetReqT {pkt: .pkt}: begin
        int_metadata$switch_id <= 'h0;
        int_metadata$insert_byte_cnt <= 'h0;
        int_metadata$insert_cnt <= 'h0;
        int_metadata$gpe_int_hdr_len8 <= 'h0;
        int_metadata$gpe_int_hdr_len <= 'h0;
        int_metadata$instruction_cnt <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_reset_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntResetRspT {pkt: pkt, int_metadata$switch_id: int_metadata$switch_id, int_metadata$gpe_int_hdr_len8: int_metadata$gpe_int_hdr_len8, int_metadata$insert_cnt: int_metadata$insert_cnt, int_metadata$gpe_int_hdr_len: int_metadata$gpe_int_hdr_len, int_metadata$insert_byte_cnt: int_metadata$insert_byte_cnt, int_metadata$instruction_cnt: int_metadata$instruction_cnt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_E_BIT ======

interface IntSetEBit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetEBit  (IntSetEBit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_header$e <- mkReg(0);
  rule int_set_e_bit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetEBitReqT {pkt: .pkt}: begin
        int_header$e <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_e_bit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetEBitRspT {pkt: pkt, int_header$e: int_header$e};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I0 ======

interface IntSetHeader0003I0;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I0  (IntSetHeader0003I0);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule int_set_header_0003_i0_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I0ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i0_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I0RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I1 ======

interface IntSetHeader0003I1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I1  (IntSetHeader0003I1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(7)) int_q_occupancy_header$q_occupancy1 <- mkReg(0);
  Reg#(Bit#(24)) int_q_occupancy_header$q_occupancy0 <- mkReg(0);
  rule int_set_header_0003_i1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I1ReqT {pkt: .pkt, intrinsic_metadata$enq_qdepth: .intrinsic_metadata$enq_qdepth}: begin
        int_q_occupancy_header$q_occupancy1 <= 'h0;
        int_q_occupancy_header$q_occupancy0 <= intrinsic_metadata$enq_qdepth;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I1RspT {pkt: pkt, int_q_occupancy_header$q_occupancy0: int_q_occupancy_header$q_occupancy0, int_q_occupancy_header$q_occupancy1: int_q_occupancy_header$q_occupancy1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I10 ======

interface IntSetHeader0003I10;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I10  (IntSetHeader0003I10);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_hop_latency_header$hop_latency <- mkReg(0);
  Reg#(Bit#(31)) int_switch_id_header$switch_id <- mkReg(0);
  rule int_set_header_0003_i10_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I10ReqT {pkt: .pkt, intrinsic_metadata$deq_timedelta: .intrinsic_metadata$deq_timedelta, int_metadata$switch_id: .int_metadata$switch_id}: begin
        int_hop_latency_header$hop_latency <= intrinsic_metadata$deq_timedelta;
        int_switch_id_header$switch_id <= int_metadata$switch_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i10_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I10RspT {pkt: pkt, int_switch_id_header$switch_id: int_switch_id_header$switch_id, int_hop_latency_header$hop_latency: int_hop_latency_header$hop_latency};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I11 ======

interface IntSetHeader0003I11;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I11  (IntSetHeader0003I11);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(7)) int_q_occupancy_header$q_occupancy1 <- mkReg(0);
  Reg#(Bit#(24)) int_q_occupancy_header$q_occupancy0 <- mkReg(0);
  Reg#(Bit#(31)) int_hop_latency_header$hop_latency <- mkReg(0);
  Reg#(Bit#(31)) int_switch_id_header$switch_id <- mkReg(0);
  rule int_set_header_0003_i11_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I11ReqT {pkt: .pkt, intrinsic_metadata$deq_timedelta: .intrinsic_metadata$deq_timedelta, intrinsic_metadata$enq_qdepth: .intrinsic_metadata$enq_qdepth, int_metadata$switch_id: .int_metadata$switch_id}: begin
        int_q_occupancy_header$q_occupancy1 <= 'h0;
        int_q_occupancy_header$q_occupancy0 <= intrinsic_metadata$enq_qdepth;
        int_hop_latency_header$hop_latency <= intrinsic_metadata$deq_timedelta;
        int_switch_id_header$switch_id <= int_metadata$switch_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i11_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I11RspT {pkt: pkt, int_switch_id_header$switch_id: int_switch_id_header$switch_id, int_q_occupancy_header$q_occupancy0: int_q_occupancy_header$q_occupancy0, int_hop_latency_header$hop_latency: int_hop_latency_header$hop_latency, int_q_occupancy_header$q_occupancy1: int_q_occupancy_header$q_occupancy1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I12 ======

interface IntSetHeader0003I12;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I12  (IntSetHeader0003I12);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(15)) int_ingress_port_id_header$ingress_port_id_1 <- mkReg(0);
  Reg#(Bit#(16)) int_ingress_port_id_header$ingress_port_id_0 <- mkReg(0);
  Reg#(Bit#(31)) int_switch_id_header$switch_id <- mkReg(0);
  rule int_set_header_0003_i12_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I12ReqT {pkt: .pkt, int_metadata$switch_id: .int_metadata$switch_id, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        int_ingress_port_id_header$ingress_port_id_1 <= 'h0;
        int_ingress_port_id_header$ingress_port_id_0 <= ingress_metadata$ifindex;
        int_switch_id_header$switch_id <= int_metadata$switch_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i12_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I12RspT {pkt: pkt, int_ingress_port_id_header$ingress_port_id_1: int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: int_ingress_port_id_header$ingress_port_id_0, int_switch_id_header$switch_id: int_switch_id_header$switch_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I13 ======

interface IntSetHeader0003I13;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I13  (IntSetHeader0003I13);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(7)) int_q_occupancy_header$q_occupancy1 <- mkReg(0);
  Reg#(Bit#(24)) int_q_occupancy_header$q_occupancy0 <- mkReg(0);
  Reg#(Bit#(15)) int_ingress_port_id_header$ingress_port_id_1 <- mkReg(0);
  Reg#(Bit#(16)) int_ingress_port_id_header$ingress_port_id_0 <- mkReg(0);
  Reg#(Bit#(31)) int_switch_id_header$switch_id <- mkReg(0);
  rule int_set_header_0003_i13_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I13ReqT {pkt: .pkt, int_metadata$switch_id: .int_metadata$switch_id, intrinsic_metadata$enq_qdepth: .intrinsic_metadata$enq_qdepth, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        int_q_occupancy_header$q_occupancy1 <= 'h0;
        int_q_occupancy_header$q_occupancy0 <= intrinsic_metadata$enq_qdepth;
        int_ingress_port_id_header$ingress_port_id_1 <= 'h0;
        int_ingress_port_id_header$ingress_port_id_0 <= ingress_metadata$ifindex;
        int_switch_id_header$switch_id <= int_metadata$switch_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i13_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I13RspT {pkt: pkt, int_ingress_port_id_header$ingress_port_id_1: int_ingress_port_id_header$ingress_port_id_1, int_q_occupancy_header$q_occupancy0: int_q_occupancy_header$q_occupancy0, int_ingress_port_id_header$ingress_port_id_0: int_ingress_port_id_header$ingress_port_id_0, int_switch_id_header$switch_id: int_switch_id_header$switch_id, int_q_occupancy_header$q_occupancy1: int_q_occupancy_header$q_occupancy1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I14 ======

interface IntSetHeader0003I14;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I14  (IntSetHeader0003I14);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_hop_latency_header$hop_latency <- mkReg(0);
  Reg#(Bit#(15)) int_ingress_port_id_header$ingress_port_id_1 <- mkReg(0);
  Reg#(Bit#(16)) int_ingress_port_id_header$ingress_port_id_0 <- mkReg(0);
  Reg#(Bit#(31)) int_switch_id_header$switch_id <- mkReg(0);
  rule int_set_header_0003_i14_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I14ReqT {pkt: .pkt, intrinsic_metadata$deq_timedelta: .intrinsic_metadata$deq_timedelta, ingress_metadata$ifindex: .ingress_metadata$ifindex, int_metadata$switch_id: .int_metadata$switch_id}: begin
        int_hop_latency_header$hop_latency <= intrinsic_metadata$deq_timedelta;
        int_ingress_port_id_header$ingress_port_id_1 <= 'h0;
        int_ingress_port_id_header$ingress_port_id_0 <= ingress_metadata$ifindex;
        int_switch_id_header$switch_id <= int_metadata$switch_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i14_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I14RspT {pkt: pkt, int_ingress_port_id_header$ingress_port_id_1: int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: int_ingress_port_id_header$ingress_port_id_0, int_switch_id_header$switch_id: int_switch_id_header$switch_id, int_hop_latency_header$hop_latency: int_hop_latency_header$hop_latency};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I15 ======

interface IntSetHeader0003I15;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I15  (IntSetHeader0003I15);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(7)) int_q_occupancy_header$q_occupancy1 <- mkReg(0);
  Reg#(Bit#(24)) int_q_occupancy_header$q_occupancy0 <- mkReg(0);
  Reg#(Bit#(31)) int_hop_latency_header$hop_latency <- mkReg(0);
  Reg#(Bit#(15)) int_ingress_port_id_header$ingress_port_id_1 <- mkReg(0);
  Reg#(Bit#(16)) int_ingress_port_id_header$ingress_port_id_0 <- mkReg(0);
  Reg#(Bit#(31)) int_switch_id_header$switch_id <- mkReg(0);
  rule int_set_header_0003_i15_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I15ReqT {pkt: .pkt, intrinsic_metadata$deq_timedelta: .intrinsic_metadata$deq_timedelta, intrinsic_metadata$enq_qdepth: .intrinsic_metadata$enq_qdepth, ingress_metadata$ifindex: .ingress_metadata$ifindex, int_metadata$switch_id: .int_metadata$switch_id}: begin
        int_q_occupancy_header$q_occupancy1 <= 'h0;
        int_q_occupancy_header$q_occupancy0 <= intrinsic_metadata$enq_qdepth;
        int_hop_latency_header$hop_latency <= intrinsic_metadata$deq_timedelta;
        int_ingress_port_id_header$ingress_port_id_1 <= 'h0;
        int_ingress_port_id_header$ingress_port_id_0 <= ingress_metadata$ifindex;
        int_switch_id_header$switch_id <= int_metadata$switch_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i15_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I15RspT {pkt: pkt, int_q_occupancy_header$q_occupancy0: int_q_occupancy_header$q_occupancy0, int_switch_id_header$switch_id: int_switch_id_header$switch_id, int_hop_latency_header$hop_latency: int_hop_latency_header$hop_latency, int_ingress_port_id_header$ingress_port_id_1: int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: int_ingress_port_id_header$ingress_port_id_0, int_q_occupancy_header$q_occupancy1: int_q_occupancy_header$q_occupancy1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I2 ======

interface IntSetHeader0003I2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I2  (IntSetHeader0003I2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_hop_latency_header$hop_latency <- mkReg(0);
  rule int_set_header_0003_i2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I2ReqT {pkt: .pkt, intrinsic_metadata$deq_timedelta: .intrinsic_metadata$deq_timedelta}: begin
        int_hop_latency_header$hop_latency <= intrinsic_metadata$deq_timedelta;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I2RspT {pkt: pkt, int_hop_latency_header$hop_latency: int_hop_latency_header$hop_latency};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I3 ======

interface IntSetHeader0003I3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I3  (IntSetHeader0003I3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(7)) int_q_occupancy_header$q_occupancy1 <- mkReg(0);
  Reg#(Bit#(24)) int_q_occupancy_header$q_occupancy0 <- mkReg(0);
  Reg#(Bit#(31)) int_hop_latency_header$hop_latency <- mkReg(0);
  rule int_set_header_0003_i3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I3ReqT {pkt: .pkt, intrinsic_metadata$deq_timedelta: .intrinsic_metadata$deq_timedelta, intrinsic_metadata$enq_qdepth: .intrinsic_metadata$enq_qdepth}: begin
        int_q_occupancy_header$q_occupancy1 <= 'h0;
        int_q_occupancy_header$q_occupancy0 <= intrinsic_metadata$enq_qdepth;
        int_hop_latency_header$hop_latency <= intrinsic_metadata$deq_timedelta;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I3RspT {pkt: pkt, int_q_occupancy_header$q_occupancy0: int_q_occupancy_header$q_occupancy0, int_hop_latency_header$hop_latency: int_hop_latency_header$hop_latency, int_q_occupancy_header$q_occupancy1: int_q_occupancy_header$q_occupancy1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I4 ======

interface IntSetHeader0003I4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I4  (IntSetHeader0003I4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(15)) int_ingress_port_id_header$ingress_port_id_1 <- mkReg(0);
  Reg#(Bit#(16)) int_ingress_port_id_header$ingress_port_id_0 <- mkReg(0);
  rule int_set_header_0003_i4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I4ReqT {pkt: .pkt, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        int_ingress_port_id_header$ingress_port_id_1 <= 'h0;
        int_ingress_port_id_header$ingress_port_id_0 <= ingress_metadata$ifindex;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I4RspT {pkt: pkt, int_ingress_port_id_header$ingress_port_id_1: int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: int_ingress_port_id_header$ingress_port_id_0};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I5 ======

interface IntSetHeader0003I5;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I5  (IntSetHeader0003I5);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(7)) int_q_occupancy_header$q_occupancy1 <- mkReg(0);
  Reg#(Bit#(24)) int_q_occupancy_header$q_occupancy0 <- mkReg(0);
  Reg#(Bit#(15)) int_ingress_port_id_header$ingress_port_id_1 <- mkReg(0);
  Reg#(Bit#(16)) int_ingress_port_id_header$ingress_port_id_0 <- mkReg(0);
  rule int_set_header_0003_i5_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I5ReqT {pkt: .pkt, intrinsic_metadata$enq_qdepth: .intrinsic_metadata$enq_qdepth, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        int_q_occupancy_header$q_occupancy1 <= 'h0;
        int_q_occupancy_header$q_occupancy0 <= intrinsic_metadata$enq_qdepth;
        int_ingress_port_id_header$ingress_port_id_1 <= 'h0;
        int_ingress_port_id_header$ingress_port_id_0 <= ingress_metadata$ifindex;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i5_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I5RspT {pkt: pkt, int_ingress_port_id_header$ingress_port_id_1: int_ingress_port_id_header$ingress_port_id_1, int_q_occupancy_header$q_occupancy0: int_q_occupancy_header$q_occupancy0, int_ingress_port_id_header$ingress_port_id_0: int_ingress_port_id_header$ingress_port_id_0, int_q_occupancy_header$q_occupancy1: int_q_occupancy_header$q_occupancy1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I6 ======

interface IntSetHeader0003I6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I6  (IntSetHeader0003I6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_hop_latency_header$hop_latency <- mkReg(0);
  Reg#(Bit#(15)) int_ingress_port_id_header$ingress_port_id_1 <- mkReg(0);
  Reg#(Bit#(16)) int_ingress_port_id_header$ingress_port_id_0 <- mkReg(0);
  rule int_set_header_0003_i6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I6ReqT {pkt: .pkt, intrinsic_metadata$deq_timedelta: .intrinsic_metadata$deq_timedelta, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        int_hop_latency_header$hop_latency <= intrinsic_metadata$deq_timedelta;
        int_ingress_port_id_header$ingress_port_id_1 <= 'h0;
        int_ingress_port_id_header$ingress_port_id_0 <= ingress_metadata$ifindex;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I6RspT {pkt: pkt, int_ingress_port_id_header$ingress_port_id_1: int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: int_ingress_port_id_header$ingress_port_id_0, int_hop_latency_header$hop_latency: int_hop_latency_header$hop_latency};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I7 ======

interface IntSetHeader0003I7;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I7  (IntSetHeader0003I7);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(7)) int_q_occupancy_header$q_occupancy1 <- mkReg(0);
  Reg#(Bit#(24)) int_q_occupancy_header$q_occupancy0 <- mkReg(0);
  Reg#(Bit#(31)) int_hop_latency_header$hop_latency <- mkReg(0);
  Reg#(Bit#(15)) int_ingress_port_id_header$ingress_port_id_1 <- mkReg(0);
  Reg#(Bit#(16)) int_ingress_port_id_header$ingress_port_id_0 <- mkReg(0);
  rule int_set_header_0003_i7_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I7ReqT {pkt: .pkt, intrinsic_metadata$deq_timedelta: .intrinsic_metadata$deq_timedelta, intrinsic_metadata$enq_qdepth: .intrinsic_metadata$enq_qdepth, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        int_q_occupancy_header$q_occupancy1 <= 'h0;
        int_q_occupancy_header$q_occupancy0 <= intrinsic_metadata$enq_qdepth;
        int_hop_latency_header$hop_latency <= intrinsic_metadata$deq_timedelta;
        int_ingress_port_id_header$ingress_port_id_1 <= 'h0;
        int_ingress_port_id_header$ingress_port_id_0 <= ingress_metadata$ifindex;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i7_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I7RspT {pkt: pkt, int_ingress_port_id_header$ingress_port_id_1: int_ingress_port_id_header$ingress_port_id_1, int_q_occupancy_header$q_occupancy0: int_q_occupancy_header$q_occupancy0, int_ingress_port_id_header$ingress_port_id_0: int_ingress_port_id_header$ingress_port_id_0, int_hop_latency_header$hop_latency: int_hop_latency_header$hop_latency, int_q_occupancy_header$q_occupancy1: int_q_occupancy_header$q_occupancy1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I8 ======

interface IntSetHeader0003I8;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I8  (IntSetHeader0003I8);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_switch_id_header$switch_id <- mkReg(0);
  rule int_set_header_0003_i8_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I8ReqT {pkt: .pkt, int_metadata$switch_id: .int_metadata$switch_id}: begin
        int_switch_id_header$switch_id <= int_metadata$switch_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i8_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I8RspT {pkt: pkt, int_switch_id_header$switch_id: int_switch_id_header$switch_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0003_I9 ======

interface IntSetHeader0003I9;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0003I9  (IntSetHeader0003I9);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(7)) int_q_occupancy_header$q_occupancy1 <- mkReg(0);
  Reg#(Bit#(24)) int_q_occupancy_header$q_occupancy0 <- mkReg(0);
  Reg#(Bit#(31)) int_switch_id_header$switch_id <- mkReg(0);
  rule int_set_header_0003_i9_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0003I9ReqT {pkt: .pkt, int_metadata$switch_id: .int_metadata$switch_id, intrinsic_metadata$enq_qdepth: .intrinsic_metadata$enq_qdepth}: begin
        int_q_occupancy_header$q_occupancy1 <= 'h0;
        int_q_occupancy_header$q_occupancy0 <= intrinsic_metadata$enq_qdepth;
        int_switch_id_header$switch_id <= int_metadata$switch_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0003_i9_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0003I9RspT {pkt: pkt, int_q_occupancy_header$q_occupancy0: int_q_occupancy_header$q_occupancy0, int_switch_id_header$switch_id: int_switch_id_header$switch_id, int_q_occupancy_header$q_occupancy1: int_q_occupancy_header$q_occupancy1};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I0 ======

interface IntSetHeader0407I0;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I0  (IntSetHeader0407I0);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule int_set_header_0407_i0_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I0ReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i0_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I0RspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I1 ======

interface IntSetHeader0407I1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I1  (IntSetHeader0407I1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_tx_utilization_header$egress_port_tx_utilization <- mkReg(0);
  rule int_set_header_0407_i1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I1ReqT {pkt: .pkt}: begin
        int_egress_port_tx_utilization_header$egress_port_tx_utilization <= 'h7fffffff;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I1RspT {pkt: pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: int_egress_port_tx_utilization_header$egress_port_tx_utilization};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I10 ======

interface IntSetHeader0407I10;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I10  (IntSetHeader0407I10);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_q_congestion_header$q_congestion <- mkReg(0);
  Reg#(Bit#(31)) int_ingress_tstamp_header$ingress_tstamp <- mkReg(0);
  rule int_set_header_0407_i10_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I10ReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp}: begin
        int_q_congestion_header$q_congestion <= 'h7fffffff;
        int_ingress_tstamp_header$ingress_tstamp <= i2e_metadata$ingress_tstamp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i10_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I10RspT {pkt: pkt, int_q_congestion_header$q_congestion: int_q_congestion_header$q_congestion, int_ingress_tstamp_header$ingress_tstamp: int_ingress_tstamp_header$ingress_tstamp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I11 ======

interface IntSetHeader0407I11;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I11  (IntSetHeader0407I11);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_tx_utilization_header$egress_port_tx_utilization <- mkReg(0);
  Reg#(Bit#(31)) int_q_congestion_header$q_congestion <- mkReg(0);
  Reg#(Bit#(31)) int_ingress_tstamp_header$ingress_tstamp <- mkReg(0);
  rule int_set_header_0407_i11_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I11ReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp}: begin
        int_egress_port_tx_utilization_header$egress_port_tx_utilization <= 'h7fffffff;
        int_q_congestion_header$q_congestion <= 'h7fffffff;
        int_ingress_tstamp_header$ingress_tstamp <= i2e_metadata$ingress_tstamp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i11_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I11RspT {pkt: pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_q_congestion_header$q_congestion: int_q_congestion_header$q_congestion, int_ingress_tstamp_header$ingress_tstamp: int_ingress_tstamp_header$ingress_tstamp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I12 ======

interface IntSetHeader0407I12;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I12  (IntSetHeader0407I12);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_id_header$egress_port_id <- mkReg(0);
  Reg#(Bit#(31)) int_ingress_tstamp_header$ingress_tstamp <- mkReg(0);
  rule int_set_header_0407_i12_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I12ReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, standard_metadata$egress_port: .standard_metadata$egress_port}: begin
        int_egress_port_id_header$egress_port_id <= standard_metadata$egress_port;
        int_ingress_tstamp_header$ingress_tstamp <= i2e_metadata$ingress_tstamp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i12_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I12RspT {pkt: pkt, int_egress_port_id_header$egress_port_id: int_egress_port_id_header$egress_port_id, int_ingress_tstamp_header$ingress_tstamp: int_ingress_tstamp_header$ingress_tstamp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I13 ======

interface IntSetHeader0407I13;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I13  (IntSetHeader0407I13);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_tx_utilization_header$egress_port_tx_utilization <- mkReg(0);
  Reg#(Bit#(31)) int_egress_port_id_header$egress_port_id <- mkReg(0);
  Reg#(Bit#(31)) int_ingress_tstamp_header$ingress_tstamp <- mkReg(0);
  rule int_set_header_0407_i13_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I13ReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, standard_metadata$egress_port: .standard_metadata$egress_port}: begin
        int_egress_port_tx_utilization_header$egress_port_tx_utilization <= 'h7fffffff;
        int_egress_port_id_header$egress_port_id <= standard_metadata$egress_port;
        int_ingress_tstamp_header$ingress_tstamp <= i2e_metadata$ingress_tstamp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i13_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I13RspT {pkt: pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_egress_port_id_header$egress_port_id: int_egress_port_id_header$egress_port_id, int_ingress_tstamp_header$ingress_tstamp: int_ingress_tstamp_header$ingress_tstamp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I14 ======

interface IntSetHeader0407I14;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I14  (IntSetHeader0407I14);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_q_congestion_header$q_congestion <- mkReg(0);
  Reg#(Bit#(31)) int_egress_port_id_header$egress_port_id <- mkReg(0);
  Reg#(Bit#(31)) int_ingress_tstamp_header$ingress_tstamp <- mkReg(0);
  rule int_set_header_0407_i14_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I14ReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, standard_metadata$egress_port: .standard_metadata$egress_port}: begin
        int_q_congestion_header$q_congestion <= 'h7fffffff;
        int_egress_port_id_header$egress_port_id <= standard_metadata$egress_port;
        int_ingress_tstamp_header$ingress_tstamp <= i2e_metadata$ingress_tstamp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i14_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I14RspT {pkt: pkt, int_q_congestion_header$q_congestion: int_q_congestion_header$q_congestion, int_egress_port_id_header$egress_port_id: int_egress_port_id_header$egress_port_id, int_ingress_tstamp_header$ingress_tstamp: int_ingress_tstamp_header$ingress_tstamp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I15 ======

interface IntSetHeader0407I15;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I15  (IntSetHeader0407I15);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_tx_utilization_header$egress_port_tx_utilization <- mkReg(0);
  Reg#(Bit#(31)) int_q_congestion_header$q_congestion <- mkReg(0);
  Reg#(Bit#(31)) int_egress_port_id_header$egress_port_id <- mkReg(0);
  Reg#(Bit#(31)) int_ingress_tstamp_header$ingress_tstamp <- mkReg(0);
  rule int_set_header_0407_i15_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I15ReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, standard_metadata$egress_port: .standard_metadata$egress_port}: begin
        int_egress_port_tx_utilization_header$egress_port_tx_utilization <= 'h7fffffff;
        int_q_congestion_header$q_congestion <= 'h7fffffff;
        int_egress_port_id_header$egress_port_id <= standard_metadata$egress_port;
        int_ingress_tstamp_header$ingress_tstamp <= i2e_metadata$ingress_tstamp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i15_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I15RspT {pkt: pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_egress_port_id_header$egress_port_id: int_egress_port_id_header$egress_port_id, int_q_congestion_header$q_congestion: int_q_congestion_header$q_congestion, int_ingress_tstamp_header$ingress_tstamp: int_ingress_tstamp_header$ingress_tstamp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I2 ======

interface IntSetHeader0407I2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I2  (IntSetHeader0407I2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_q_congestion_header$q_congestion <- mkReg(0);
  rule int_set_header_0407_i2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I2ReqT {pkt: .pkt}: begin
        int_q_congestion_header$q_congestion <= 'h7fffffff;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I2RspT {pkt: pkt, int_q_congestion_header$q_congestion: int_q_congestion_header$q_congestion};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I3 ======

interface IntSetHeader0407I3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I3  (IntSetHeader0407I3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_tx_utilization_header$egress_port_tx_utilization <- mkReg(0);
  Reg#(Bit#(31)) int_q_congestion_header$q_congestion <- mkReg(0);
  rule int_set_header_0407_i3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I3ReqT {pkt: .pkt}: begin
        int_egress_port_tx_utilization_header$egress_port_tx_utilization <= 'h7fffffff;
        int_q_congestion_header$q_congestion <= 'h7fffffff;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I3RspT {pkt: pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_q_congestion_header$q_congestion: int_q_congestion_header$q_congestion};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I4 ======

interface IntSetHeader0407I4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I4  (IntSetHeader0407I4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_id_header$egress_port_id <- mkReg(0);
  rule int_set_header_0407_i4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I4ReqT {pkt: .pkt, standard_metadata$egress_port: .standard_metadata$egress_port}: begin
        int_egress_port_id_header$egress_port_id <= standard_metadata$egress_port;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I4RspT {pkt: pkt, int_egress_port_id_header$egress_port_id: int_egress_port_id_header$egress_port_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I5 ======

interface IntSetHeader0407I5;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I5  (IntSetHeader0407I5);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_tx_utilization_header$egress_port_tx_utilization <- mkReg(0);
  Reg#(Bit#(31)) int_egress_port_id_header$egress_port_id <- mkReg(0);
  rule int_set_header_0407_i5_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I5ReqT {pkt: .pkt, standard_metadata$egress_port: .standard_metadata$egress_port}: begin
        int_egress_port_tx_utilization_header$egress_port_tx_utilization <= 'h7fffffff;
        int_egress_port_id_header$egress_port_id <= standard_metadata$egress_port;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i5_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I5RspT {pkt: pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_egress_port_id_header$egress_port_id: int_egress_port_id_header$egress_port_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I6 ======

interface IntSetHeader0407I6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I6  (IntSetHeader0407I6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_q_congestion_header$q_congestion <- mkReg(0);
  Reg#(Bit#(31)) int_egress_port_id_header$egress_port_id <- mkReg(0);
  rule int_set_header_0407_i6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I6ReqT {pkt: .pkt, standard_metadata$egress_port: .standard_metadata$egress_port}: begin
        int_q_congestion_header$q_congestion <= 'h7fffffff;
        int_egress_port_id_header$egress_port_id <= standard_metadata$egress_port;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I6RspT {pkt: pkt, int_q_congestion_header$q_congestion: int_q_congestion_header$q_congestion, int_egress_port_id_header$egress_port_id: int_egress_port_id_header$egress_port_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I7 ======

interface IntSetHeader0407I7;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I7  (IntSetHeader0407I7);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_tx_utilization_header$egress_port_tx_utilization <- mkReg(0);
  Reg#(Bit#(31)) int_q_congestion_header$q_congestion <- mkReg(0);
  Reg#(Bit#(31)) int_egress_port_id_header$egress_port_id <- mkReg(0);
  rule int_set_header_0407_i7_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I7ReqT {pkt: .pkt, standard_metadata$egress_port: .standard_metadata$egress_port}: begin
        int_egress_port_tx_utilization_header$egress_port_tx_utilization <= 'h7fffffff;
        int_q_congestion_header$q_congestion <= 'h7fffffff;
        int_egress_port_id_header$egress_port_id <= standard_metadata$egress_port;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i7_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I7RspT {pkt: pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_egress_port_id_header$egress_port_id: int_egress_port_id_header$egress_port_id, int_q_congestion_header$q_congestion: int_q_congestion_header$q_congestion};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I8 ======

interface IntSetHeader0407I8;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I8  (IntSetHeader0407I8);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_ingress_tstamp_header$ingress_tstamp <- mkReg(0);
  rule int_set_header_0407_i8_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I8ReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp}: begin
        int_ingress_tstamp_header$ingress_tstamp <= i2e_metadata$ingress_tstamp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i8_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I8RspT {pkt: pkt, int_ingress_tstamp_header$ingress_tstamp: int_ingress_tstamp_header$ingress_tstamp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0407_I9 ======

interface IntSetHeader0407I9;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0407I9  (IntSetHeader0407I9);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(31)) int_egress_port_tx_utilization_header$egress_port_tx_utilization <- mkReg(0);
  Reg#(Bit#(31)) int_ingress_tstamp_header$ingress_tstamp <- mkReg(0);
  rule int_set_header_0407_i9_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0407I9ReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp}: begin
        int_egress_port_tx_utilization_header$egress_port_tx_utilization <= 'h7fffffff;
        int_ingress_tstamp_header$ingress_tstamp <= i2e_metadata$ingress_tstamp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0407_i9_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0407I9RspT {pkt: pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_ingress_tstamp_header$ingress_tstamp: int_ingress_tstamp_header$ingress_tstamp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_0_BOS ======

interface IntSetHeader0Bos;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader0Bos  (IntSetHeader0Bos);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_switch_id_header$bos <- mkReg(0);
  rule int_set_header_0_bos_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader0BosReqT {pkt: .pkt}: begin
        int_switch_id_header$bos <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_0_bos_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader0BosRspT {pkt: pkt, int_switch_id_header$bos: int_switch_id_header$bos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_1_BOS ======

interface IntSetHeader1Bos;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader1Bos  (IntSetHeader1Bos);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_ingress_port_id_header$bos <- mkReg(0);
  rule int_set_header_1_bos_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader1BosReqT {pkt: .pkt}: begin
        int_ingress_port_id_header$bos <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_1_bos_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader1BosRspT {pkt: pkt, int_ingress_port_id_header$bos: int_ingress_port_id_header$bos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_2_BOS ======

interface IntSetHeader2Bos;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader2Bos  (IntSetHeader2Bos);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_hop_latency_header$bos <- mkReg(0);
  rule int_set_header_2_bos_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader2BosReqT {pkt: .pkt}: begin
        int_hop_latency_header$bos <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_2_bos_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader2BosRspT {pkt: pkt, int_hop_latency_header$bos: int_hop_latency_header$bos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_3_BOS ======

interface IntSetHeader3Bos;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader3Bos  (IntSetHeader3Bos);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_q_occupancy_header$bos <- mkReg(0);
  rule int_set_header_3_bos_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader3BosReqT {pkt: .pkt}: begin
        int_q_occupancy_header$bos <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_3_bos_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader3BosRspT {pkt: pkt, int_q_occupancy_header$bos: int_q_occupancy_header$bos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_4_BOS ======

interface IntSetHeader4Bos;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader4Bos  (IntSetHeader4Bos);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_ingress_tstamp_header$bos <- mkReg(0);
  rule int_set_header_4_bos_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader4BosReqT {pkt: .pkt}: begin
        int_ingress_tstamp_header$bos <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_4_bos_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader4BosRspT {pkt: pkt, int_ingress_tstamp_header$bos: int_ingress_tstamp_header$bos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_5_BOS ======

interface IntSetHeader5Bos;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader5Bos  (IntSetHeader5Bos);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_egress_port_id_header$bos <- mkReg(0);
  rule int_set_header_5_bos_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader5BosReqT {pkt: .pkt}: begin
        int_egress_port_id_header$bos <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_5_bos_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader5BosRspT {pkt: pkt, int_egress_port_id_header$bos: int_egress_port_id_header$bos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_6_BOS ======

interface IntSetHeader6Bos;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader6Bos  (IntSetHeader6Bos);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_q_congestion_header$bos <- mkReg(0);
  rule int_set_header_6_bos_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader6BosReqT {pkt: .pkt}: begin
        int_q_congestion_header$bos <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_6_bos_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader6BosRspT {pkt: pkt, int_q_congestion_header$bos: int_q_congestion_header$bos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_HEADER_7_BOS ======

interface IntSetHeader7Bos;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetHeader7Bos  (IntSetHeader7Bos);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_egress_port_tx_utilization_header$bos <- mkReg(0);
  rule int_set_header_7_bos_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetHeader7BosReqT {pkt: .pkt}: begin
        int_egress_port_tx_utilization_header$bos <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_header_7_bos_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetHeader7BosRspT {pkt: pkt, int_egress_port_tx_utilization_header$bos: int_egress_port_tx_utilization_header$bos};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_NO_SRC ======

interface IntSetNoSrc;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetNoSrc  (IntSetNoSrc);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_metadata_i2e$source <- mkReg(0);
  rule int_set_no_src_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetNoSrcReqT {pkt: .pkt}: begin
        int_metadata_i2e$source <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_no_src_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetNoSrcRspT {pkt: pkt, int_metadata_i2e$source: int_metadata_i2e$source};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SET_SRC ======

interface IntSetSrc;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSetSrc  (IntSetSrc);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_metadata_i2e$source <- mkReg(0);
  rule int_set_src_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSetSrcReqT {pkt: .pkt}: begin
        int_metadata_i2e$source <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_set_src_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSetSrcRspT {pkt: pkt, int_metadata_i2e$source: int_metadata_i2e$source};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SINK_GPE ======

interface IntSinkGpe;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSinkGpe  (IntSinkGpe);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) int_metadata_i2e$sink <- mkReg(0);
  Reg#(Bit#(16)) i2e_metadata$mirror_session_id <- mkReg(0);
  rule int_sink_gpe_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSinkGpeReqT {pkt: .pkt, runtime_mirror_id: .runtime_mirror_id}: begin
        int_metadata_i2e$sink <= 'h1;
        i2e_metadata$mirror_session_id <= runtime_mirror_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_sink_gpe_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSinkGpeRspT {pkt: pkt, i2e_metadata$mirror_session_id: i2e_metadata$mirror_session_id, int_metadata_i2e$sink: int_metadata_i2e$sink};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SINK_UPDATE_VXLAN_GPE_V4 ======

interface IntSinkUpdateVxlanGpeV4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSinkUpdateVxlanGpeV4  (IntSinkUpdateVxlanGpeV4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) vxlan_gpe$next_proto <- mkReg(0);
  rule int_sink_update_vxlan_gpe_v4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSinkUpdateVxlanGpeV4ReqT {pkt: .pkt, vxlan_gpe_int_header$next_proto: .vxlan_gpe_int_header$next_proto}: begin
        vxlan_gpe$next_proto <= vxlan_gpe_int_header$next_proto;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_sink_update_vxlan_gpe_v4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSinkUpdateVxlanGpeV4RspT {pkt: pkt, vxlan_gpe$next_proto: vxlan_gpe$next_proto};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_SRC ======

interface IntSrc;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntSrc  (IntSrc);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) int_metadata$insert_cnt <- mkReg(0);
  Reg#(Bit#(32)) int_metadata$switch_id <- mkReg(0);
  Reg#(Bit#(16)) int_metadata$insert_byte_cnt <- mkReg(0);
  Reg#(Bit#(8)) int_metadata$gpe_int_hdr_len8 <- mkReg(0);
  Reg#(Bit#(2)) int_header$ver <- mkReg(0);
  Reg#(Bit#(2)) int_header$rep <- mkReg(0);
  Reg#(Bit#(1)) int_header$c <- mkReg(0);
  Reg#(Bit#(1)) int_header$e <- mkReg(0);
  Reg#(Bit#(5)) int_header$rsvd1 <- mkReg(0);
  Reg#(Bit#(5)) int_header$ins_cnt <- mkReg(0);
  Reg#(Bit#(8)) int_header$max_hop_cnt <- mkReg(0);
  Reg#(Bit#(8)) int_header$total_hop_cnt <- mkReg(0);
  Reg#(Bit#(4)) int_header$instruction_mask_0003 <- mkReg(0);
  Reg#(Bit#(4)) int_header$instruction_mask_0407 <- mkReg(0);
  Reg#(Bit#(4)) int_header$instruction_mask_0811 <- mkReg(0);
  Reg#(Bit#(4)) int_header$instruction_mask_1215 <- mkReg(0);
  Reg#(Bit#(16)) int_header$rsvd2 <- mkReg(0);
  rule int_src_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntSrcReqT {pkt: .pkt, runtime_total_words: .runtime_total_words, runtime_switch_id: .runtime_switch_id, runtime_ins_mask0003: .runtime_ins_mask0003, runtime_ins_byte_cnt: .runtime_ins_byte_cnt, runtime_ins_cnt: .runtime_ins_cnt, runtime_hop_cnt: .runtime_hop_cnt, runtime_ins_mask0407: .runtime_ins_mask0407}: begin
        int_metadata$insert_cnt <= runtime_hop_cnt;
        int_metadata$switch_id <= runtime_switch_id;
        int_metadata$insert_byte_cnt <= runtime_ins_byte_cnt;
        int_metadata$gpe_int_hdr_len8 <= runtime_total_words;
        int_header$ver <= 'h0;
        int_header$rep <= 'h0;
        int_header$c <= 'h0;
        int_header$e <= 'h0;
        int_header$rsvd1 <= 'h0;
        int_header$ins_cnt <= runtime_ins_cnt;
        int_header$max_hop_cnt <= runtime_hop_cnt;
        int_header$total_hop_cnt <= 'h0;
        int_header$instruction_mask_0003 <= runtime_ins_mask0003;
        int_header$instruction_mask_0407 <= runtime_ins_mask0407;
        int_header$instruction_mask_0811 <= 'h0;
        int_header$instruction_mask_1215 <= 'h0;
        int_header$rsvd2 <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_src_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntSrcRspT {pkt: pkt, int_metadata$gpe_int_hdr_len8: int_metadata$gpe_int_hdr_len8, int_header$rsvd2: int_header$rsvd2, int_header$ins_cnt: int_header$ins_cnt, int_header$instruction_mask_0407: int_header$instruction_mask_0407, int_header$total_hop_cnt: int_header$total_hop_cnt, int_header$instruction_mask_1215: int_header$instruction_mask_1215, int_header$rsvd1: int_header$rsvd1, int_header$e: int_header$e, int_header$instruction_mask_0811: int_header$instruction_mask_0811, int_metadata$switch_id: int_metadata$switch_id, int_header$rep: int_header$rep, int_header$ver: int_header$ver, int_header$max_hop_cnt: int_header$max_hop_cnt, int_header$instruction_mask_0003: int_header$instruction_mask_0003, int_metadata$insert_cnt: int_metadata$insert_cnt, int_header$c: int_header$c, int_metadata$insert_byte_cnt: int_metadata$insert_byte_cnt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_TRANSIT ======

interface IntTransit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntTransit  (IntTransit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(32)) int_metadata$switch_id <- mkReg(0);
  Reg#(Bit#(8)) int_metadata$gpe_int_hdr_len8 <- mkReg(0);
  rule int_transit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntTransitReqT {pkt: .pkt, int_header$ins_cnt: .int_header$ins_cnt, runtime_switch_id: .runtime_switch_id}: begin
        int_metadata$switch_id <= runtime_switch_id;
        int_metadata$gpe_int_hdr_len8 <= int_header$ins_cnt;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_transit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntTransitRspT {pkt: pkt, int_metadata$switch_id: int_metadata$switch_id, int_metadata$gpe_int_hdr_len8: int_metadata$gpe_int_hdr_len8};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_UPDATE_TOTAL_HOP_CNT ======

interface IntUpdateTotalHopCnt;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntUpdateTotalHopCnt  (IntUpdateTotalHopCnt);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule int_update_total_hop_cnt_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntUpdateTotalHopCntReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_update_total_hop_cnt_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntUpdateTotalHopCntRspT {pkt: pkt, int_header$total_hop_cnt: int_header$total_hop_cnt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== INT_UPDATE_VXLAN_GPE_IPV4 ======

interface IntUpdateVxlanGpeIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIntUpdateVxlanGpeIpv4  (IntUpdateVxlanGpeIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule int_update_vxlan_gpe_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IntUpdateVxlanGpeIpv4ReqT {pkt: .pkt, int_metadata$gpe_int_hdr_len8: .int_metadata$gpe_int_hdr_len8, int_metadata$insert_byte_cnt: .int_metadata$insert_byte_cnt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule int_update_vxlan_gpe_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IntUpdateVxlanGpeIpv4RspT {pkt: pkt, vxlan_gpe_int_header$len: vxlan_gpe_int_header$len, udp$length_: udp$length_, ipv4$totalLen: ipv4$totalLen};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPSG_MISS ======

interface IpsgMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpsgMiss  (IpsgMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) security_metadata$ipsg_check_fail <- mkReg(0);
  rule ipsg_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged IpsgMissReqT {pkt: .pkt}: begin
        security_metadata$ipsg_check_fail <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipsg_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged IpsgMissRspT {pkt: pkt, security_metadata$ipsg_check_fail: security_metadata$ipsg_check_fail};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_ERSPAN_T3_REWRITE ======

interface Ipv4ErspanT3Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4ErspanT3Rewrite  (Ipv4ErspanT3Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) gre$C <- mkReg(0);
  Reg#(Bit#(1)) gre$R <- mkReg(0);
  Reg#(Bit#(1)) gre$K <- mkReg(0);
  Reg#(Bit#(1)) gre$S <- mkReg(0);
  Reg#(Bit#(1)) gre$s <- mkReg(0);
  Reg#(Bit#(3)) gre$recurse <- mkReg(0);
  Reg#(Bit#(5)) gre$flags <- mkReg(0);
  Reg#(Bit#(3)) gre$ver <- mkReg(0);
  Reg#(Bit#(16)) gre$proto <- mkReg(0);
  Reg#(Bit#(32)) erspan_t3_header$timestamp <- mkReg(0);
  Reg#(Bit#(10)) erspan_t3_header$span_id <- mkReg(0);
  Reg#(Bit#(4)) erspan_t3_header$version <- mkReg(0);
  Reg#(Bit#(32)) erspan_t3_header$sgt_other <- mkReg(0);
  Reg#(Bit#(8)) ipv4$protocol <- mkReg(0);
  Reg#(Bit#(8)) ipv4$ttl <- mkReg(0);
  Reg#(Bit#(4)) ipv4$version <- mkReg(0);
  Reg#(Bit#(4)) ipv4$ihl <- mkReg(0);
  Reg#(Bit#(16)) ipv4$identification <- mkReg(0);
  rule ipv4_erspan_t3_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4ErspanT3RewriteReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id}: begin
        gre$C <= 'h0;
        gre$R <= 'h0;
        gre$K <= 'h0;
        gre$S <= 'h0;
        gre$s <= 'h0;
        gre$recurse <= 'h0;
        gre$flags <= 'h0;
        gre$ver <= 'h0;
        gre$proto <= 'h22eb;
        erspan_t3_header$timestamp <= i2e_metadata$ingress_tstamp;
        erspan_t3_header$span_id <= i2e_metadata$mirror_session_id;
        erspan_t3_header$version <= 'h2;
        erspan_t3_header$sgt_other <= 'h0;
        ipv4$protocol <= 'h2f;
        ipv4$ttl <= 'h40;
        ipv4$version <= 'h4;
        ipv4$ihl <= 'h5;
        ipv4$identification <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_erspan_t3_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4ErspanT3RewriteRspT {pkt: pkt, gre$S: gre$S, ipv4$identification: ipv4$identification, gre$s: gre$s, ipv4$version: ipv4$version, ipv4$ihl: ipv4$ihl, gre$proto: gre$proto, ipv4$ttl: ipv4$ttl, gre$ver: gre$ver, erspan_t3_header$timestamp: erspan_t3_header$timestamp, gre$C: gre$C, gre$recurse: gre$recurse, erspan_t3_header$span_id: erspan_t3_header$span_id, gre$K: gre$K, erspan_t3_header$version: erspan_t3_header$version, gre$flags: gre$flags, erspan_t3_header$sgt_other: erspan_t3_header$sgt_other, ipv4$protocol: ipv4$protocol, gre$R: gre$R};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_GENV_REWRITE ======

interface Ipv4GenvRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4GenvRewrite  (Ipv4GenvRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) udp$srcPort <- mkReg(0);
  Reg#(Bit#(16)) udp$dstPort <- mkReg(0);
  Reg#(Bit#(16)) udp$checksum <- mkReg(0);
  Reg#(Bit#(2)) genv$ver <- mkReg(0);
  Reg#(Bit#(1)) genv$oam <- mkReg(0);
  Reg#(Bit#(1)) genv$critical <- mkReg(0);
  Reg#(Bit#(6)) genv$optLen <- mkReg(0);
  Reg#(Bit#(16)) genv$protoType <- mkReg(0);
  Reg#(Bit#(24)) genv$vni <- mkReg(0);
  Reg#(Bit#(6)) genv$reserved <- mkReg(0);
  Reg#(Bit#(8)) genv$reserved2 <- mkReg(0);
  Reg#(Bit#(8)) ipv4$protocol <- mkReg(0);
  Reg#(Bit#(8)) ipv4$ttl <- mkReg(0);
  Reg#(Bit#(4)) ipv4$version <- mkReg(0);
  Reg#(Bit#(4)) ipv4$ihl <- mkReg(0);
  Reg#(Bit#(16)) ipv4$identification <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv4_genv_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4GenvRewriteReqT {pkt: .pkt, hash_metadata$entropy_hash: .hash_metadata$entropy_hash, tunnel_metadata$vnid: .tunnel_metadata$vnid}: begin
        udp$srcPort <= hash_metadata$entropy_hash;
        udp$dstPort <= 'h17c1;
        udp$checksum <= 'h0;
        genv$ver <= 'h0;
        genv$oam <= 'h0;
        genv$critical <= 'h0;
        genv$optLen <= 'h0;
        genv$protoType <= 'h6558;
        genv$vni <= tunnel_metadata$vnid;
        genv$reserved <= 'h0;
        genv$reserved2 <= 'h0;
        ipv4$protocol <= 'h11;
        ipv4$ttl <= 'h40;
        ipv4$version <= 'h4;
        ipv4$ihl <= 'h5;
        ipv4$identification <= 'h0;
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_genv_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4GenvRewriteRspT {pkt: pkt, genv$vni: genv$vni, ipv4$identification: ipv4$identification, udp$checksum: udp$checksum, ipv4$version: ipv4$version, ipv4$ihl: ipv4$ihl, genv$optLen: genv$optLen, ipv4$ttl: ipv4$ttl, genv$oam: genv$oam, genv$reserved2: genv$reserved2, genv$critical: genv$critical, udp$srcPort: udp$srcPort, genv$protoType: genv$protoType, genv$ver: genv$ver, udp$dstPort: udp$dstPort, ethernet$etherType: ethernet$etherType, ipv4$protocol: ipv4$protocol, genv$reserved: genv$reserved};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_GRE_REWRITE ======

interface Ipv4GreRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4GreRewrite  (Ipv4GreRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) gre$proto <- mkReg(0);
  Reg#(Bit#(8)) ipv4$protocol <- mkReg(0);
  Reg#(Bit#(8)) ipv4$ttl <- mkReg(0);
  Reg#(Bit#(4)) ipv4$version <- mkReg(0);
  Reg#(Bit#(4)) ipv4$ihl <- mkReg(0);
  Reg#(Bit#(16)) ipv4$identification <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv4_gre_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4GreRewriteReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        gre$proto <= ethernet$etherType;
        ipv4$protocol <= 'h2f;
        ipv4$ttl <= 'h40;
        ipv4$version <= 'h4;
        ipv4$ihl <= 'h5;
        ipv4$identification <= 'h0;
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_gre_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4GreRewriteRspT {pkt: pkt, ipv4$protocol: ipv4$protocol, ipv4$ihl: ipv4$ihl, gre$proto: gre$proto, ipv4$ttl: ipv4$ttl, ipv4$identification: ipv4$identification, ethernet$etherType: ethernet$etherType, ipv4$version: ipv4$version};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_IP_REWRITE ======

interface Ipv4IpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4IpRewrite  (Ipv4IpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) ipv4$protocol <- mkReg(0);
  Reg#(Bit#(8)) ipv4$ttl <- mkReg(0);
  Reg#(Bit#(4)) ipv4$version <- mkReg(0);
  Reg#(Bit#(4)) ipv4$ihl <- mkReg(0);
  Reg#(Bit#(16)) ipv4$identification <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv4_ip_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4IpRewriteReqT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto}: begin
        ipv4$protocol <= tunnel_metadata$inner_ip_proto;
        ipv4$ttl <= 'h40;
        ipv4$version <= 'h4;
        ipv4$ihl <= 'h5;
        ipv4$identification <= 'h0;
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_ip_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4IpRewriteRspT {pkt: pkt, ipv4$protocol: ipv4$protocol, ipv4$ihl: ipv4$ihl, ipv4$ttl: ipv4$ttl, ipv4$identification: ipv4$identification, ethernet$etherType: ethernet$etherType, ipv4$version: ipv4$version};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_MTU_CHECK ======

interface Ipv4MtuCheck;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4MtuCheck  (Ipv4MtuCheck);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule ipv4_mtu_check_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4MtuCheckReqT {pkt: .pkt, runtime_l3_mtu: .runtime_l3_mtu}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_mtu_check_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4MtuCheckRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_MULTICAST_REWRITE ======

interface Ipv4MulticastRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4MulticastRewrite  (Ipv4MulticastRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule ipv4_multicast_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4MulticastRewriteReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_multicast_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4MulticastRewriteRspT {pkt: pkt, ipv4$ttl: ipv4$ttl};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_NVGRE_REWRITE ======

interface Ipv4NvgreRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4NvgreRewrite  (Ipv4NvgreRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) gre$proto <- mkReg(0);
  Reg#(Bit#(3)) gre$recurse <- mkReg(0);
  Reg#(Bit#(5)) gre$flags <- mkReg(0);
  Reg#(Bit#(3)) gre$ver <- mkReg(0);
  Reg#(Bit#(1)) gre$R <- mkReg(0);
  Reg#(Bit#(1)) gre$K <- mkReg(0);
  Reg#(Bit#(1)) gre$C <- mkReg(0);
  Reg#(Bit#(1)) gre$S <- mkReg(0);
  Reg#(Bit#(1)) gre$s <- mkReg(0);
  Reg#(Bit#(24)) nvgre$tni <- mkReg(0);
  Reg#(Bit#(8)) nvgre$flow_id <- mkReg(0);
  Reg#(Bit#(8)) ipv4$protocol <- mkReg(0);
  Reg#(Bit#(8)) ipv4$ttl <- mkReg(0);
  Reg#(Bit#(4)) ipv4$version <- mkReg(0);
  Reg#(Bit#(4)) ipv4$ihl <- mkReg(0);
  Reg#(Bit#(16)) ipv4$identification <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv4_nvgre_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4NvgreRewriteReqT {pkt: .pkt, tunnel_metadata$vnid: .tunnel_metadata$vnid}: begin
        gre$proto <= 'h6558;
        gre$recurse <= 'h0;
        gre$flags <= 'h0;
        gre$ver <= 'h0;
        gre$R <= 'h0;
        gre$K <= 'h1;
        gre$C <= 'h0;
        gre$S <= 'h0;
        gre$s <= 'h0;
        nvgre$tni <= tunnel_metadata$vnid;
        nvgre$flow_id <= type$value;
        ipv4$protocol <= 'h2f;
        ipv4$ttl <= 'h40;
        ipv4$version <= 'h4;
        ipv4$ihl <= 'h5;
        ipv4$identification <= 'h0;
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_nvgre_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4NvgreRewriteRspT {pkt: pkt, gre$s: gre$s, ipv4$identification: ipv4$identification, gre$R: gre$R, nvgre$flow_id: nvgre$flow_id, ipv4$ihl: ipv4$ihl, gre$proto: gre$proto, ipv4$ttl: ipv4$ttl, gre$ver: gre$ver, gre$S: gre$S, gre$C: gre$C, gre$recurse: gre$recurse, nvgre$tni: nvgre$tni, gre$K: gre$K, gre$flags: gre$flags, ethernet$etherType: ethernet$etherType, ipv4$protocol: ipv4$protocol, ipv4$version: ipv4$version};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_OVER_FABRIC ======

interface Ipv4OverFabric;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4OverFabric  (Ipv4OverFabric);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(32)) ipv4_metadata$lkp_ipv4_sa <- mkReg(0);
  Reg#(Bit#(32)) ipv4_metadata$lkp_ipv4_da <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_proto <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$lkp_l4_sport <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$lkp_l4_dport <- mkReg(0);
  rule ipv4_over_fabric_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4OverFabricReqT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, ipv4$srcAddr: .ipv4$srcAddr, ipv4$dstAddr: .ipv4$dstAddr, l3_metadata$lkp_outer_l4_dport: .l3_metadata$lkp_outer_l4_dport, ipv4$protocol: .ipv4$protocol, l3_metadata$lkp_outer_l4_sport: .l3_metadata$lkp_outer_l4_sport}: begin
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        ipv4_metadata$lkp_ipv4_sa <= ipv4$srcAddr;
        ipv4_metadata$lkp_ipv4_da <= ipv4$dstAddr;
        l3_metadata$lkp_ip_proto <= ipv4$protocol;
        l3_metadata$lkp_l4_sport <= l3_metadata$lkp_outer_l4_sport;
        l3_metadata$lkp_l4_dport <= l3_metadata$lkp_outer_l4_dport;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_over_fabric_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4OverFabricRspT {pkt: pkt, ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da, ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa, l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_sport: l3_metadata$lkp_l4_sport, l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_TUNNEL_LOOKUP_MISS ======

interface Ipv4TunnelLookupMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4TunnelLookupMiss  (Ipv4TunnelLookupMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(32)) ipv4_metadata$lkp_ipv4_sa <- mkReg(0);
  Reg#(Bit#(32)) ipv4_metadata$lkp_ipv4_da <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_proto <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_ttl <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$lkp_l4_sport <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$lkp_l4_dport <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  rule ipv4_tunnel_lookup_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4TunnelLookupMissReqT {pkt: .pkt, l3_metadata$lkp_outer_l4_dport: .l3_metadata$lkp_outer_l4_dport, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, ipv4$srcAddr: .ipv4$srcAddr, ipv4$dstAddr: .ipv4$dstAddr, ipv4$ttl: .ipv4$ttl, ipv4$protocol: .ipv4$protocol, l3_metadata$lkp_outer_l4_sport: .l3_metadata$lkp_outer_l4_sport}: begin
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        ipv4_metadata$lkp_ipv4_sa <= ipv4$srcAddr;
        ipv4_metadata$lkp_ipv4_da <= ipv4$dstAddr;
        l3_metadata$lkp_ip_proto <= ipv4$protocol;
        l3_metadata$lkp_ip_ttl <= ipv4$ttl;
        l3_metadata$lkp_l4_sport <= l3_metadata$lkp_outer_l4_sport;
        l3_metadata$lkp_l4_dport <= l3_metadata$lkp_outer_l4_dport;
        intrinsic_metadata$mcast_grp <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_tunnel_lookup_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4TunnelLookupMissRspT {pkt: pkt, l3_metadata$lkp_ip_ttl: l3_metadata$lkp_ip_ttl, ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da, ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_sport: l3_metadata$lkp_l4_sport, l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_UNICAST_REWRITE ======

interface Ipv4UnicastRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4UnicastRewrite  (Ipv4UnicastRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) ethernet$dstAddr <- mkReg(0);
  rule ipv4_unicast_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4UnicastRewriteReqT {pkt: .pkt, egress_metadata$mac_da: .egress_metadata$mac_da}: begin
        ethernet$dstAddr <= egress_metadata$mac_da;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_unicast_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4UnicastRewriteRspT {pkt: pkt, ipv4$ttl: ipv4$ttl, ethernet$dstAddr: ethernet$dstAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_URPF_HIT ======

interface Ipv4UrpfHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4UrpfHit  (Ipv4UrpfHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$urpf_hit <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$urpf_bd_group <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$urpf_mode <- mkReg(0);
  rule ipv4_urpf_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4UrpfHitReqT {pkt: .pkt, ipv4_metadata$ipv4_urpf_mode: .ipv4_metadata$ipv4_urpf_mode, runtime_urpf_bd_group: .runtime_urpf_bd_group}: begin
        l3_metadata$urpf_hit <= 'h1;
        l3_metadata$urpf_bd_group <= runtime_urpf_bd_group;
        l3_metadata$urpf_mode <= ipv4_metadata$ipv4_urpf_mode;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_urpf_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4UrpfHitRspT {pkt: pkt, l3_metadata$urpf_bd_group: l3_metadata$urpf_bd_group, l3_metadata$urpf_hit: l3_metadata$urpf_hit, l3_metadata$urpf_mode: l3_metadata$urpf_mode};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV4_VXLAN_REWRITE ======

interface Ipv4VxlanRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv4VxlanRewrite  (Ipv4VxlanRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) udp$srcPort <- mkReg(0);
  Reg#(Bit#(16)) udp$dstPort <- mkReg(0);
  Reg#(Bit#(16)) udp$checksum <- mkReg(0);
  Reg#(Bit#(None)) vxlan$flags <- mkReg(0);
  Reg#(Bit#(None)) vxlan$reserved <- mkReg(0);
  Reg#(Bit#(None)) vxlan$vni <- mkReg(0);
  Reg#(Bit#(None)) vxlan$reserved2 <- mkReg(0);
  Reg#(Bit#(8)) ipv4$protocol <- mkReg(0);
  Reg#(Bit#(8)) ipv4$ttl <- mkReg(0);
  Reg#(Bit#(4)) ipv4$version <- mkReg(0);
  Reg#(Bit#(4)) ipv4$ihl <- mkReg(0);
  Reg#(Bit#(16)) ipv4$identification <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv4_vxlan_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv4VxlanRewriteReqT {pkt: .pkt, hash_metadata$entropy_hash: .hash_metadata$entropy_hash, tunnel_metadata$vnid: .tunnel_metadata$vnid}: begin
        udp$srcPort <= hash_metadata$entropy_hash;
        udp$dstPort <= 'h12b5;
        udp$checksum <= 'h0;
        vxlan$flags <= 'h8;
        vxlan$reserved <= 'h0;
        vxlan$vni <= tunnel_metadata$vnid;
        vxlan$reserved2 <= 'h0;
        ipv4$protocol <= 'h11;
        ipv4$ttl <= 'h40;
        ipv4$version <= 'h4;
        ipv4$ihl <= 'h5;
        ipv4$identification <= 'h0;
        ethernet$etherType <= 'h800;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv4_vxlan_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv4VxlanRewriteRspT {pkt: pkt, ipv4$identification: ipv4$identification, udp$checksum: udp$checksum, vxlan$vni: vxlan$vni, ipv4$ihl: ipv4$ihl, vxlan$flags: vxlan$flags, ipv4$ttl: ipv4$ttl, ipv4$protocol: ipv4$protocol, vxlan$reserved2: vxlan$reserved2, udp$srcPort: udp$srcPort, vxlan$reserved: vxlan$reserved, udp$dstPort: udp$dstPort, ethernet$etherType: ethernet$etherType, ipv4$version: ipv4$version};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_ERSPAN_T3_REWRITE ======

interface Ipv6ErspanT3Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6ErspanT3Rewrite  (Ipv6ErspanT3Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) gre$C <- mkReg(0);
  Reg#(Bit#(1)) gre$R <- mkReg(0);
  Reg#(Bit#(1)) gre$K <- mkReg(0);
  Reg#(Bit#(1)) gre$S <- mkReg(0);
  Reg#(Bit#(1)) gre$s <- mkReg(0);
  Reg#(Bit#(3)) gre$recurse <- mkReg(0);
  Reg#(Bit#(5)) gre$flags <- mkReg(0);
  Reg#(Bit#(3)) gre$ver <- mkReg(0);
  Reg#(Bit#(16)) gre$proto <- mkReg(0);
  Reg#(Bit#(32)) erspan_t3_header$timestamp <- mkReg(0);
  Reg#(Bit#(10)) erspan_t3_header$span_id <- mkReg(0);
  Reg#(Bit#(4)) erspan_t3_header$version <- mkReg(0);
  Reg#(Bit#(32)) erspan_t3_header$sgt_other <- mkReg(0);
  Reg#(Bit#(4)) ipv6$version <- mkReg(0);
  Reg#(Bit#(8)) ipv6$nextHdr <- mkReg(0);
  Reg#(Bit#(8)) ipv6$hopLimit <- mkReg(0);
  Reg#(Bit#(8)) ipv6$trafficClass <- mkReg(0);
  Reg#(Bit#(20)) ipv6$flowLabel <- mkReg(0);
  rule ipv6_erspan_t3_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6ErspanT3RewriteReqT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id}: begin
        gre$C <= 'h0;
        gre$R <= 'h0;
        gre$K <= 'h0;
        gre$S <= 'h0;
        gre$s <= 'h0;
        gre$recurse <= 'h0;
        gre$flags <= 'h0;
        gre$ver <= 'h0;
        gre$proto <= 'h22eb;
        erspan_t3_header$timestamp <= i2e_metadata$ingress_tstamp;
        erspan_t3_header$span_id <= i2e_metadata$mirror_session_id;
        erspan_t3_header$version <= 'h2;
        erspan_t3_header$sgt_other <= 'h0;
        ipv6$version <= 'h6;
        ipv6$nextHdr <= 'h2f;
        ipv6$hopLimit <= 'h40;
        ipv6$trafficClass <= 'h0;
        ipv6$flowLabel <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_erspan_t3_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6ErspanT3RewriteRspT {pkt: pkt, ipv6$version: ipv6$version, gre$S: gre$S, ipv6$trafficClass: ipv6$trafficClass, gre$s: gre$s, ipv6$hopLimit: ipv6$hopLimit, ipv6$flowLabel: ipv6$flowLabel, gre$proto: gre$proto, gre$ver: gre$ver, erspan_t3_header$timestamp: erspan_t3_header$timestamp, gre$C: gre$C, gre$recurse: gre$recurse, ipv6$nextHdr: ipv6$nextHdr, erspan_t3_header$span_id: erspan_t3_header$span_id, gre$K: gre$K, erspan_t3_header$version: erspan_t3_header$version, gre$flags: gre$flags, erspan_t3_header$sgt_other: erspan_t3_header$sgt_other, gre$R: gre$R};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_GENV_REWRITE ======

interface Ipv6GenvRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6GenvRewrite  (Ipv6GenvRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) udp$srcPort <- mkReg(0);
  Reg#(Bit#(16)) udp$dstPort <- mkReg(0);
  Reg#(Bit#(16)) udp$checksum <- mkReg(0);
  Reg#(Bit#(2)) genv$ver <- mkReg(0);
  Reg#(Bit#(1)) genv$oam <- mkReg(0);
  Reg#(Bit#(1)) genv$critical <- mkReg(0);
  Reg#(Bit#(6)) genv$optLen <- mkReg(0);
  Reg#(Bit#(16)) genv$protoType <- mkReg(0);
  Reg#(Bit#(24)) genv$vni <- mkReg(0);
  Reg#(Bit#(6)) genv$reserved <- mkReg(0);
  Reg#(Bit#(8)) genv$reserved2 <- mkReg(0);
  Reg#(Bit#(4)) ipv6$version <- mkReg(0);
  Reg#(Bit#(8)) ipv6$nextHdr <- mkReg(0);
  Reg#(Bit#(8)) ipv6$hopLimit <- mkReg(0);
  Reg#(Bit#(8)) ipv6$trafficClass <- mkReg(0);
  Reg#(Bit#(20)) ipv6$flowLabel <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv6_genv_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6GenvRewriteReqT {pkt: .pkt, hash_metadata$entropy_hash: .hash_metadata$entropy_hash, tunnel_metadata$vnid: .tunnel_metadata$vnid}: begin
        udp$srcPort <= hash_metadata$entropy_hash;
        udp$dstPort <= 'h17c1;
        udp$checksum <= 'h0;
        genv$ver <= 'h0;
        genv$oam <= 'h0;
        genv$critical <= 'h0;
        genv$optLen <= 'h0;
        genv$protoType <= 'h6558;
        genv$vni <= tunnel_metadata$vnid;
        genv$reserved <= 'h0;
        genv$reserved2 <= 'h0;
        ipv6$version <= 'h6;
        ipv6$nextHdr <= 'h11;
        ipv6$hopLimit <= 'h40;
        ipv6$trafficClass <= 'h0;
        ipv6$flowLabel <= 'h0;
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_genv_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6GenvRewriteRspT {pkt: pkt, genv$vni: genv$vni, ipv6$trafficClass: ipv6$trafficClass, udp$checksum: udp$checksum, ipv6$version: ipv6$version, genv$optLen: genv$optLen, ipv6$nextHdr: ipv6$nextHdr, genv$oam: genv$oam, genv$reserved2: genv$reserved2, ethernet$etherType: ethernet$etherType, genv$critical: genv$critical, udp$srcPort: udp$srcPort, ipv6$flowLabel: ipv6$flowLabel, genv$protoType: genv$protoType, genv$ver: genv$ver, udp$dstPort: udp$dstPort, ipv6$hopLimit: ipv6$hopLimit, genv$reserved: genv$reserved};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_GRE_REWRITE ======

interface Ipv6GreRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6GreRewrite  (Ipv6GreRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) gre$proto <- mkReg(0);
  Reg#(Bit#(4)) ipv6$version <- mkReg(0);
  Reg#(Bit#(8)) ipv6$nextHdr <- mkReg(0);
  Reg#(Bit#(8)) ipv6$hopLimit <- mkReg(0);
  Reg#(Bit#(8)) ipv6$trafficClass <- mkReg(0);
  Reg#(Bit#(20)) ipv6$flowLabel <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv6_gre_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6GreRewriteReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        gre$proto <= ethernet$etherType;
        ipv6$version <= 'h6;
        ipv6$nextHdr <= 'h2f;
        ipv6$hopLimit <= 'h40;
        ipv6$trafficClass <= 'h0;
        ipv6$flowLabel <= 'h0;
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_gre_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6GreRewriteRspT {pkt: pkt, ipv6$version: ipv6$version, ipv6$flowLabel: ipv6$flowLabel, gre$proto: gre$proto, ipv6$hopLimit: ipv6$hopLimit, ipv6$trafficClass: ipv6$trafficClass, ipv6$nextHdr: ipv6$nextHdr, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_IP_REWRITE ======

interface Ipv6IpRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6IpRewrite  (Ipv6IpRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(4)) ipv6$version <- mkReg(0);
  Reg#(Bit#(8)) ipv6$nextHdr <- mkReg(0);
  Reg#(Bit#(8)) ipv6$hopLimit <- mkReg(0);
  Reg#(Bit#(8)) ipv6$trafficClass <- mkReg(0);
  Reg#(Bit#(20)) ipv6$flowLabel <- mkReg(0);
  Reg#(Bit#(16)) ipv6$payloadLen <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv6_ip_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6IpRewriteReqT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: .egress_metadata$payload_length}: begin
        ipv6$version <= 'h6;
        ipv6$nextHdr <= tunnel_metadata$inner_ip_proto;
        ipv6$hopLimit <= 'h40;
        ipv6$trafficClass <= 'h0;
        ipv6$flowLabel <= 'h0;
        ipv6$payloadLen <= egress_metadata$payload_length;
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_ip_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6IpRewriteRspT {pkt: pkt, ipv6$version: ipv6$version, ipv6$payloadLen: ipv6$payloadLen, ipv6$flowLabel: ipv6$flowLabel, ipv6$hopLimit: ipv6$hopLimit, ipv6$trafficClass: ipv6$trafficClass, ipv6$nextHdr: ipv6$nextHdr, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_MTU_CHECK ======

interface Ipv6MtuCheck;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6MtuCheck  (Ipv6MtuCheck);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule ipv6_mtu_check_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6MtuCheckReqT {pkt: .pkt, runtime_l3_mtu: .runtime_l3_mtu}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_mtu_check_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6MtuCheckRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_MULTICAST_REWRITE ======

interface Ipv6MulticastRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6MulticastRewrite  (Ipv6MulticastRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule ipv6_multicast_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6MulticastRewriteReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_multicast_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6MulticastRewriteRspT {pkt: pkt, ipv6$hopLimit: ipv6$hopLimit};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_NVGRE_REWRITE ======

interface Ipv6NvgreRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6NvgreRewrite  (Ipv6NvgreRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) gre$proto <- mkReg(0);
  Reg#(Bit#(3)) gre$recurse <- mkReg(0);
  Reg#(Bit#(5)) gre$flags <- mkReg(0);
  Reg#(Bit#(3)) gre$ver <- mkReg(0);
  Reg#(Bit#(1)) gre$R <- mkReg(0);
  Reg#(Bit#(1)) gre$K <- mkReg(0);
  Reg#(Bit#(1)) gre$C <- mkReg(0);
  Reg#(Bit#(1)) gre$S <- mkReg(0);
  Reg#(Bit#(1)) gre$s <- mkReg(0);
  Reg#(Bit#(24)) nvgre$tni <- mkReg(0);
  Reg#(Bit#(8)) nvgre$flow_id <- mkReg(0);
  Reg#(Bit#(4)) ipv6$version <- mkReg(0);
  Reg#(Bit#(8)) ipv6$nextHdr <- mkReg(0);
  Reg#(Bit#(8)) ipv6$hopLimit <- mkReg(0);
  Reg#(Bit#(8)) ipv6$trafficClass <- mkReg(0);
  Reg#(Bit#(20)) ipv6$flowLabel <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv6_nvgre_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6NvgreRewriteReqT {pkt: .pkt, tunnel_metadata$vnid: .tunnel_metadata$vnid}: begin
        gre$proto <= 'h6558;
        gre$recurse <= 'h0;
        gre$flags <= 'h0;
        gre$ver <= 'h0;
        gre$R <= 'h0;
        gre$K <= 'h1;
        gre$C <= 'h0;
        gre$S <= 'h0;
        gre$s <= 'h0;
        nvgre$tni <= tunnel_metadata$vnid;
        nvgre$flow_id <= type$value;
        ipv6$version <= 'h6;
        ipv6$nextHdr <= 'h2f;
        ipv6$hopLimit <= 'h40;
        ipv6$trafficClass <= 'h0;
        ipv6$flowLabel <= 'h0;
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_nvgre_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6NvgreRewriteRspT {pkt: pkt, ipv6$version: ipv6$version, gre$s: gre$s, gre$R: gre$R, nvgre$flow_id: nvgre$flow_id, gre$proto: gre$proto, gre$ver: gre$ver, gre$S: gre$S, ethernet$etherType: ethernet$etherType, gre$C: gre$C, gre$recurse: gre$recurse, nvgre$tni: nvgre$tni, ipv6$nextHdr: ipv6$nextHdr, ipv6$flowLabel: ipv6$flowLabel, gre$K: gre$K, ipv6$trafficClass: ipv6$trafficClass, gre$flags: gre$flags, ipv6$hopLimit: ipv6$hopLimit};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_OVER_FABRIC ======

interface Ipv6OverFabric;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6OverFabric  (Ipv6OverFabric);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(128)) ipv6_metadata$lkp_ipv6_sa <- mkReg(0);
  Reg#(Bit#(128)) ipv6_metadata$lkp_ipv6_da <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_proto <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$lkp_l4_sport <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$lkp_l4_dport <- mkReg(0);
  rule ipv6_over_fabric_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6OverFabricReqT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, ipv6$srcAddr: .ipv6$srcAddr, l3_metadata$lkp_outer_l4_dport: .l3_metadata$lkp_outer_l4_dport, ipv6$dstAddr: .ipv6$dstAddr, ipv6$nextHdr: .ipv6$nextHdr, l3_metadata$lkp_outer_l4_sport: .l3_metadata$lkp_outer_l4_sport}: begin
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        ipv6_metadata$lkp_ipv6_sa <= ipv6$srcAddr;
        ipv6_metadata$lkp_ipv6_da <= ipv6$dstAddr;
        l3_metadata$lkp_ip_proto <= ipv6$nextHdr;
        l3_metadata$lkp_l4_sport <= l3_metadata$lkp_outer_l4_sport;
        l3_metadata$lkp_l4_dport <= l3_metadata$lkp_outer_l4_dport;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_over_fabric_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6OverFabricRspT {pkt: pkt, ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa, ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da, l3_metadata$lkp_l4_sport: l3_metadata$lkp_l4_sport, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport, l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_TUNNEL_LOOKUP_MISS ======

interface Ipv6TunnelLookupMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6TunnelLookupMiss  (Ipv6TunnelLookupMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(128)) ipv6_metadata$lkp_ipv6_sa <- mkReg(0);
  Reg#(Bit#(128)) ipv6_metadata$lkp_ipv6_da <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_proto <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_ttl <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$lkp_l4_sport <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$lkp_l4_dport <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  rule ipv6_tunnel_lookup_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6TunnelLookupMissReqT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, ipv6$srcAddr: .ipv6$srcAddr, l3_metadata$lkp_outer_l4_dport: .l3_metadata$lkp_outer_l4_dport, ipv6$dstAddr: .ipv6$dstAddr, ipv6$hopLimit: .ipv6$hopLimit, ipv6$nextHdr: .ipv6$nextHdr, l3_metadata$lkp_outer_l4_sport: .l3_metadata$lkp_outer_l4_sport}: begin
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        ipv6_metadata$lkp_ipv6_sa <= ipv6$srcAddr;
        ipv6_metadata$lkp_ipv6_da <= ipv6$dstAddr;
        l3_metadata$lkp_ip_proto <= ipv6$nextHdr;
        l3_metadata$lkp_ip_ttl <= ipv6$hopLimit;
        l3_metadata$lkp_l4_sport <= l3_metadata$lkp_outer_l4_sport;
        l3_metadata$lkp_l4_dport <= l3_metadata$lkp_outer_l4_dport;
        intrinsic_metadata$mcast_grp <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_tunnel_lookup_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6TunnelLookupMissRspT {pkt: pkt, ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa, ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da, l3_metadata$lkp_l4_sport: l3_metadata$lkp_l4_sport, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, l3_metadata$lkp_ip_ttl: l3_metadata$lkp_ip_ttl, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport, l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_UNICAST_REWRITE ======

interface Ipv6UnicastRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6UnicastRewrite  (Ipv6UnicastRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) ethernet$dstAddr <- mkReg(0);
  rule ipv6_unicast_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6UnicastRewriteReqT {pkt: .pkt, egress_metadata$mac_da: .egress_metadata$mac_da}: begin
        ethernet$dstAddr <= egress_metadata$mac_da;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_unicast_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6UnicastRewriteRspT {pkt: pkt, ipv6$hopLimit: ipv6$hopLimit, ethernet$dstAddr: ethernet$dstAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_URPF_HIT ======

interface Ipv6UrpfHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6UrpfHit  (Ipv6UrpfHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$urpf_hit <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$urpf_bd_group <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$urpf_mode <- mkReg(0);
  rule ipv6_urpf_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6UrpfHitReqT {pkt: .pkt, ipv6_metadata$ipv6_urpf_mode: .ipv6_metadata$ipv6_urpf_mode, runtime_urpf_bd_group: .runtime_urpf_bd_group}: begin
        l3_metadata$urpf_hit <= 'h1;
        l3_metadata$urpf_bd_group <= runtime_urpf_bd_group;
        l3_metadata$urpf_mode <= ipv6_metadata$ipv6_urpf_mode;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_urpf_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6UrpfHitRspT {pkt: pkt, l3_metadata$urpf_bd_group: l3_metadata$urpf_bd_group, l3_metadata$urpf_hit: l3_metadata$urpf_hit, l3_metadata$urpf_mode: l3_metadata$urpf_mode};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== IPV6_VXLAN_REWRITE ======

interface Ipv6VxlanRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkIpv6VxlanRewrite  (Ipv6VxlanRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) udp$srcPort <- mkReg(0);
  Reg#(Bit#(16)) udp$dstPort <- mkReg(0);
  Reg#(Bit#(16)) udp$checksum <- mkReg(0);
  Reg#(Bit#(None)) vxlan$flags <- mkReg(0);
  Reg#(Bit#(None)) vxlan$reserved <- mkReg(0);
  Reg#(Bit#(None)) vxlan$vni <- mkReg(0);
  Reg#(Bit#(None)) vxlan$reserved2 <- mkReg(0);
  Reg#(Bit#(4)) ipv6$version <- mkReg(0);
  Reg#(Bit#(8)) ipv6$nextHdr <- mkReg(0);
  Reg#(Bit#(8)) ipv6$hopLimit <- mkReg(0);
  Reg#(Bit#(8)) ipv6$trafficClass <- mkReg(0);
  Reg#(Bit#(20)) ipv6$flowLabel <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule ipv6_vxlan_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged Ipv6VxlanRewriteReqT {pkt: .pkt, hash_metadata$entropy_hash: .hash_metadata$entropy_hash, tunnel_metadata$vnid: .tunnel_metadata$vnid}: begin
        udp$srcPort <= hash_metadata$entropy_hash;
        udp$dstPort <= 'h12b5;
        udp$checksum <= 'h0;
        vxlan$flags <= 'h8;
        vxlan$reserved <= 'h0;
        vxlan$vni <= tunnel_metadata$vnid;
        vxlan$reserved2 <= 'h0;
        ipv6$version <= 'h6;
        ipv6$nextHdr <= 'h11;
        ipv6$hopLimit <= 'h40;
        ipv6$trafficClass <= 'h0;
        ipv6$flowLabel <= 'h0;
        ethernet$etherType <= 'h86dd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule ipv6_vxlan_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged Ipv6VxlanRewriteRspT {pkt: pkt, ipv6$version: ipv6$version, udp$checksum: udp$checksum, vxlan$vni: vxlan$vni, vxlan$flags: vxlan$flags, ipv6$nextHdr: ipv6$nextHdr, vxlan$reserved2: vxlan$reserved2, udp$srcPort: udp$srcPort, ipv6$flowLabel: ipv6$flowLabel, vxlan$reserved: vxlan$reserved, ipv6$hopLimit: ipv6$hopLimit, ipv6$trafficClass: ipv6$trafficClass, udp$dstPort: udp$dstPort, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MALFORMED_OUTER_ETHERNET_PACKET ======

interface MalformedOuterEthernetPacket;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMalformedOuterEthernetPacket  (MalformedOuterEthernetPacket);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) ingress_metadata$drop_flag <- mkReg(0);
  Reg#(Bit#(8)) ingress_metadata$drop_reason <- mkReg(0);
  rule malformed_outer_ethernet_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MalformedOuterEthernetPacketReqT {pkt: .pkt, runtime_drop_reason: .runtime_drop_reason}: begin
        ingress_metadata$drop_flag <= 'h1;
        ingress_metadata$drop_reason <= runtime_drop_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule malformed_outer_ethernet_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MalformedOuterEthernetPacketRspT {pkt: pkt, ingress_metadata$drop_reason: ingress_metadata$drop_reason, ingress_metadata$drop_flag: ingress_metadata$drop_flag};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== METER_DENY ======

interface MeterDeny;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMeterDeny  (MeterDeny);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule meter_deny_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MeterDenyReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule meter_deny_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MeterDenyRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== METER_PERMIT ======

interface MeterPermit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMeterPermit  (MeterPermit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule meter_permit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MeterPermitReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule meter_permit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MeterPermitRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MPLS_ETHERNET_PUSH1_REWRITE ======

interface MplsEthernetPush1Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMplsEthernetPush1Rewrite  (MplsEthernetPush1Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule mpls_ethernet_push1_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MplsEthernetPush1RewriteReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h8847;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule mpls_ethernet_push1_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MplsEthernetPush1RewriteRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MPLS_ETHERNET_PUSH2_REWRITE ======

interface MplsEthernetPush2Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMplsEthernetPush2Rewrite  (MplsEthernetPush2Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule mpls_ethernet_push2_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MplsEthernetPush2RewriteReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h8847;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule mpls_ethernet_push2_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MplsEthernetPush2RewriteRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MPLS_ETHERNET_PUSH3_REWRITE ======

interface MplsEthernetPush3Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMplsEthernetPush3Rewrite  (MplsEthernetPush3Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule mpls_ethernet_push3_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MplsEthernetPush3RewriteReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h8847;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule mpls_ethernet_push3_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MplsEthernetPush3RewriteRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MPLS_IP_PUSH1_REWRITE ======

interface MplsIpPush1Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMplsIpPush1Rewrite  (MplsIpPush1Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule mpls_ip_push1_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MplsIpPush1RewriteReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h8847;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule mpls_ip_push1_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MplsIpPush1RewriteRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MPLS_IP_PUSH2_REWRITE ======

interface MplsIpPush2Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMplsIpPush2Rewrite  (MplsIpPush2Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule mpls_ip_push2_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MplsIpPush2RewriteReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h8847;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule mpls_ip_push2_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MplsIpPush2RewriteRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MPLS_IP_PUSH3_REWRITE ======

interface MplsIpPush3Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMplsIpPush3Rewrite  (MplsIpPush3Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule mpls_ip_push3_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MplsIpPush3RewriteReqT {pkt: .pkt}: begin
        ethernet$etherType <= 'h8847;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule mpls_ip_push3_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MplsIpPush3RewriteRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MPLS_REWRITE ======

interface MplsRewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMplsRewrite  (MplsRewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) ethernet$dstAddr <- mkReg(0);
  rule mpls_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MplsRewriteReqT {pkt: .pkt, egress_metadata$mac_da: .egress_metadata$mac_da}: begin
        ethernet$dstAddr <= egress_metadata$mac_da;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule mpls_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MplsRewriteRspT {pkt: pkt, ethernet$dstAddr: ethernet$dstAddr, mpls0$ttl: mpls0$ttl};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MTU_MISS ======

interface MtuMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMtuMiss  (MtuMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) l3_metadata$l3_mtu_check <- mkReg(0);
  rule mtu_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MtuMissReqT {pkt: .pkt}: begin
        l3_metadata$l3_mtu_check <= 'hffff;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule mtu_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MtuMissRspT {pkt: pkt, l3_metadata$l3_mtu_check: l3_metadata$l3_mtu_check};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MULTICAST_BRIDGE_S_G_HIT ======

interface MulticastBridgeSGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMulticastBridgeSGHit  (MulticastBridgeSGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) multicast_metadata$multicast_bridge_mc_index <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$mcast_bridge_hit <- mkReg(0);
  rule multicast_bridge_s_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MulticastBridgeSGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index}: begin
        multicast_metadata$multicast_bridge_mc_index <= runtime_mc_index;
        multicast_metadata$mcast_bridge_hit <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule multicast_bridge_s_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MulticastBridgeSGHitRspT {pkt: pkt, multicast_metadata$mcast_bridge_hit: multicast_metadata$mcast_bridge_hit, multicast_metadata$multicast_bridge_mc_index: multicast_metadata$multicast_bridge_mc_index};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MULTICAST_BRIDGE_STAR_G_HIT ======

interface MulticastBridgeStarGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMulticastBridgeStarGHit  (MulticastBridgeStarGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) multicast_metadata$multicast_bridge_mc_index <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$mcast_bridge_hit <- mkReg(0);
  rule multicast_bridge_star_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MulticastBridgeStarGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index}: begin
        multicast_metadata$multicast_bridge_mc_index <= runtime_mc_index;
        multicast_metadata$mcast_bridge_hit <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule multicast_bridge_star_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MulticastBridgeStarGHitRspT {pkt: pkt, multicast_metadata$mcast_bridge_hit: multicast_metadata$mcast_bridge_hit, multicast_metadata$multicast_bridge_mc_index: multicast_metadata$multicast_bridge_mc_index};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MULTICAST_ROUTE_BIDIR_STAR_G_HIT ======

interface MulticastRouteBidirStarGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMulticastRouteBidirStarGHit  (MulticastRouteBidirStarGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) multicast_metadata$mcast_mode <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$multicast_route_mc_index <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$mcast_route_hit <- mkReg(0);
  rule multicast_route_bidir_star_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MulticastRouteBidirStarGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index, runtime_mcast_rpf_group: .runtime_mcast_rpf_group}: begin
        multicast_metadata$mcast_mode <= 'h2;
        multicast_metadata$multicast_route_mc_index <= runtime_mc_index;
        multicast_metadata$mcast_route_hit <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule multicast_route_bidir_star_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MulticastRouteBidirStarGHitRspT {pkt: pkt, multicast_metadata$mcast_route_hit: multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: multicast_metadata$mcast_mode};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MULTICAST_ROUTE_S_G_HIT ======

interface MulticastRouteSGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMulticastRouteSGHit  (MulticastRouteSGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) multicast_metadata$multicast_route_mc_index <- mkReg(0);
  Reg#(Bit#(2)) multicast_metadata$mcast_mode <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$mcast_route_hit <- mkReg(0);
  rule multicast_route_s_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MulticastRouteSGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index, runtime_mcast_rpf_group: .runtime_mcast_rpf_group}: begin
        multicast_metadata$multicast_route_mc_index <= runtime_mc_index;
        multicast_metadata$mcast_mode <= 'h1;
        multicast_metadata$mcast_route_hit <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule multicast_route_s_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MulticastRouteSGHitRspT {pkt: pkt, multicast_metadata$mcast_route_hit: multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: multicast_metadata$mcast_mode};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MULTICAST_ROUTE_SM_STAR_G_HIT ======

interface MulticastRouteSmStarGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMulticastRouteSmStarGHit  (MulticastRouteSmStarGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) multicast_metadata$mcast_mode <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$multicast_route_mc_index <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$mcast_route_hit <- mkReg(0);
  rule multicast_route_sm_star_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MulticastRouteSmStarGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index, runtime_mcast_rpf_group: .runtime_mcast_rpf_group}: begin
        multicast_metadata$mcast_mode <= 'h1;
        multicast_metadata$multicast_route_mc_index <= runtime_mc_index;
        multicast_metadata$mcast_route_hit <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule multicast_route_sm_star_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MulticastRouteSmStarGHitRspT {pkt: pkt, multicast_metadata$mcast_route_hit: multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: multicast_metadata$mcast_mode};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== MULTICAST_ROUTE_STAR_G_MISS ======

interface MulticastRouteStarGMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkMulticastRouteStarGMiss  (MulticastRouteStarGMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$l3_copy <- mkReg(0);
  rule multicast_route_star_g_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged MulticastRouteStarGMissReqT {pkt: .pkt}: begin
        l3_metadata$l3_copy <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule multicast_route_star_g_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged MulticastRouteStarGMissRspT {pkt: pkt, l3_metadata$l3_copy: l3_metadata$l3_copy};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== NEGATIVE_MIRROR ======

interface NegativeMirror;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkNegativeMirror  (NegativeMirror);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule negative_mirror_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged NegativeMirrorReqT {pkt: .pkt, runtime_session_id: .runtime_session_id}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule negative_mirror_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged NegativeMirrorRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== NON_IP_OVER_FABRIC ======

interface NonIpOverFabric;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkNonIpOverFabric  (NonIpOverFabric);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule non_ip_over_fabric_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged NonIpOverFabricReqT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, ethernet$etherType: .ethernet$etherType}: begin
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        l2_metadata$lkp_mac_type <= ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule non_ip_over_fabric_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged NonIpOverFabricRspT {pkt: pkt, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== NON_IP_TUNNEL_LOOKUP_MISS ======

interface NonIpTunnelLookupMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkNonIpTunnelLookupMiss  (NonIpTunnelLookupMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  rule non_ip_tunnel_lookup_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged NonIpTunnelLookupMissReqT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr}: begin
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        intrinsic_metadata$mcast_grp <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule non_ip_tunnel_lookup_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged NonIpTunnelLookupMissRspT {pkt: pkt, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== NOP ======

interface Nop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkNop  (Nop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule nop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged NopReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule nop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged NopRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== ON_MISS ======

interface OnMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkOnMiss  (OnMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule on_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged OnMissReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule on_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged OnMissRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== OUTER_MULTICAST_BRIDGE_S_G_HIT ======

interface OuterMulticastBridgeSGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkOuterMulticastBridgeSGHit  (OuterMulticastBridgeSGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule outer_multicast_bridge_s_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged OuterMulticastBridgeSGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index}: begin
        intrinsic_metadata$mcast_grp <= runtime_mc_index;
        tunnel_metadata$tunnel_terminate <= 'h1;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule outer_multicast_bridge_s_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged OuterMulticastBridgeSGHitRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== OUTER_MULTICAST_BRIDGE_STAR_G_HIT ======

interface OuterMulticastBridgeStarGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkOuterMulticastBridgeStarGHit  (OuterMulticastBridgeStarGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule outer_multicast_bridge_star_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged OuterMulticastBridgeStarGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index}: begin
        intrinsic_metadata$mcast_grp <= runtime_mc_index;
        tunnel_metadata$tunnel_terminate <= 'h1;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule outer_multicast_bridge_star_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged OuterMulticastBridgeStarGHitRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== OUTER_MULTICAST_ROUTE_BIDIR_STAR_G_HIT ======

interface OuterMulticastRouteBidirStarGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkOuterMulticastRouteBidirStarGHit  (OuterMulticastRouteBidirStarGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) multicast_metadata$outer_mcast_mode <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$outer_mcast_route_hit <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule outer_multicast_route_bidir_star_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged OuterMulticastRouteBidirStarGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index, runtime_mcast_rpf_group: .runtime_mcast_rpf_group}: begin
        multicast_metadata$outer_mcast_mode <= 'h2;
        intrinsic_metadata$mcast_grp <= runtime_mc_index;
        multicast_metadata$outer_mcast_route_hit <= 'h1;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule outer_multicast_route_bidir_star_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged OuterMulticastRouteBidirStarGHitRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: multicast_metadata$outer_mcast_route_hit, multicast_metadata$outer_mcast_mode: multicast_metadata$outer_mcast_mode, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== OUTER_MULTICAST_ROUTE_S_G_HIT ======

interface OuterMulticastRouteSGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkOuterMulticastRouteSGHit  (OuterMulticastRouteSGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$outer_mcast_route_hit <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule outer_multicast_route_s_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged OuterMulticastRouteSGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index, runtime_mcast_rpf_group: .runtime_mcast_rpf_group}: begin
        intrinsic_metadata$mcast_grp <= runtime_mc_index;
        multicast_metadata$outer_mcast_route_hit <= 'h1;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule outer_multicast_route_s_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged OuterMulticastRouteSGHitRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: multicast_metadata$outer_mcast_route_hit, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== OUTER_MULTICAST_ROUTE_SM_STAR_G_HIT ======

interface OuterMulticastRouteSmStarGHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkOuterMulticastRouteSmStarGHit  (OuterMulticastRouteSmStarGHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) multicast_metadata$outer_mcast_mode <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$outer_mcast_route_hit <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule outer_multicast_route_sm_star_g_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged OuterMulticastRouteSmStarGHitReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index, runtime_mcast_rpf_group: .runtime_mcast_rpf_group}: begin
        multicast_metadata$outer_mcast_mode <= 'h1;
        intrinsic_metadata$mcast_grp <= runtime_mc_index;
        multicast_metadata$outer_mcast_route_hit <= 'h1;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule outer_multicast_route_sm_star_g_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged OuterMulticastRouteSmStarGHitRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: multicast_metadata$outer_mcast_route_hit, multicast_metadata$outer_mcast_mode: multicast_metadata$outer_mcast_mode, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== OUTER_REPLICA_FROM_RID ======

interface OuterReplicaFromRid;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkOuterReplicaFromRid  (OuterReplicaFromRid);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$replica <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$inner_replica <- mkReg(0);
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  Reg#(Bit#(4)) tunnel_metadata$egress_header_count <- mkReg(0);
  rule outer_replica_from_rid_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged OuterReplicaFromRidReqT {pkt: .pkt, l3_metadata$outer_routed: .l3_metadata$outer_routed, runtime_tunnel_index: .runtime_tunnel_index, runtime_tunnel_type: .runtime_tunnel_type, runtime_bd: .runtime_bd, runtime_header_count: .runtime_header_count}: begin
        egress_metadata$bd <= runtime_bd;
        multicast_metadata$replica <= 'h1;
        multicast_metadata$inner_replica <= 'h0;
        egress_metadata$routed <= l3_metadata$outer_routed;
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        tunnel_metadata$egress_tunnel_type <= runtime_tunnel_type;
        tunnel_metadata$egress_header_count <= runtime_header_count;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule outer_replica_from_rid_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged OuterReplicaFromRidRspT {pkt: pkt, multicast_metadata$replica: multicast_metadata$replica, multicast_metadata$inner_replica: multicast_metadata$inner_replica, tunnel_metadata$egress_header_count: tunnel_metadata$egress_header_count, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type, egress_metadata$bd: egress_metadata$bd, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index, egress_metadata$routed: egress_metadata$routed};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== OUTER_RMAC_HIT ======

interface OuterRmacHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkOuterRmacHit  (OuterRmacHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$rmac_hit <- mkReg(0);
  rule outer_rmac_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged OuterRmacHitReqT {pkt: .pkt}: begin
        l3_metadata$rmac_hit <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule outer_rmac_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged OuterRmacHitRspT {pkt: pkt, l3_metadata$rmac_hit: l3_metadata$rmac_hit};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== PORT_VLAN_MAPPING_MISS ======

interface PortVlanMappingMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkPortVlanMappingMiss  (PortVlanMappingMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l2_metadata$port_vlan_mapping_miss <- mkReg(0);
  rule port_vlan_mapping_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged PortVlanMappingMissReqT {pkt: .pkt}: begin
        l2_metadata$port_vlan_mapping_miss <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule port_vlan_mapping_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged PortVlanMappingMissRspT {pkt: pkt, l2_metadata$port_vlan_mapping_miss: l2_metadata$port_vlan_mapping_miss};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== RACL_DENY ======

interface RaclDeny;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRaclDeny  (RaclDeny);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) acl_metadata$racl_deny <- mkReg(0);
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_copy <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule racl_deny_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RaclDenyReqT {pkt: .pkt, runtime_acl_copy: .runtime_acl_copy, runtime_acl_copy_reason: .runtime_acl_copy_reason, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        acl_metadata$racl_deny <= 'h1;
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        acl_metadata$acl_copy <= runtime_acl_copy;
        fabric_metadata$reason_code <= runtime_acl_copy_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule racl_deny_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RaclDenyRspT {pkt: pkt, acl_metadata$racl_deny: acl_metadata$racl_deny, acl_metadata$acl_copy: acl_metadata$acl_copy, fabric_metadata$reason_code: fabric_metadata$reason_code, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== RACL_PERMIT ======

interface RaclPermit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRaclPermit  (RaclPermit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_copy <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule racl_permit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RaclPermitReqT {pkt: .pkt, runtime_acl_copy: .runtime_acl_copy, runtime_acl_copy_reason: .runtime_acl_copy_reason, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        acl_metadata$acl_copy <= runtime_acl_copy;
        fabric_metadata$reason_code <= runtime_acl_copy_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule racl_permit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RaclPermitRspT {pkt: pkt, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index, acl_metadata$acl_copy: acl_metadata$acl_copy, fabric_metadata$reason_code: fabric_metadata$reason_code};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== RACL_REDIRECT_ECMP ======

interface RaclRedirectEcmp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRaclRedirectEcmp  (RaclRedirectEcmp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) acl_metadata$racl_redirect <- mkReg(0);
  Reg#(Bit#(16)) acl_metadata$racl_nexthop <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$racl_nexthop_type <- mkReg(0);
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_copy <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule racl_redirect_ecmp_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RaclRedirectEcmpReqT {pkt: .pkt, runtime_acl_copy_reason: .runtime_acl_copy_reason, runtime_acl_copy: .runtime_acl_copy, runtime_ecmp_index: .runtime_ecmp_index, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        acl_metadata$racl_redirect <= 'h1;
        acl_metadata$racl_nexthop <= runtime_ecmp_index;
        acl_metadata$racl_nexthop_type <= 'h1;
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        acl_metadata$acl_copy <= runtime_acl_copy;
        fabric_metadata$reason_code <= runtime_acl_copy_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule racl_redirect_ecmp_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RaclRedirectEcmpRspT {pkt: pkt, acl_metadata$racl_nexthop: acl_metadata$racl_nexthop, acl_metadata$acl_copy: acl_metadata$acl_copy, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index, acl_metadata$racl_redirect: acl_metadata$racl_redirect, fabric_metadata$reason_code: fabric_metadata$reason_code, acl_metadata$racl_nexthop_type: acl_metadata$racl_nexthop_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== RACL_REDIRECT_NEXTHOP ======

interface RaclRedirectNexthop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRaclRedirectNexthop  (RaclRedirectNexthop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) acl_metadata$racl_redirect <- mkReg(0);
  Reg#(Bit#(16)) acl_metadata$racl_nexthop <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$racl_nexthop_type <- mkReg(0);
  Reg#(Bit#(14)) acl_metadata$acl_stats_index <- mkReg(0);
  Reg#(Bit#(1)) acl_metadata$acl_copy <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  rule racl_redirect_nexthop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RaclRedirectNexthopReqT {pkt: .pkt, runtime_acl_copy_reason: .runtime_acl_copy_reason, runtime_acl_copy: .runtime_acl_copy, runtime_nexthop_index: .runtime_nexthop_index, runtime_acl_stats_index: .runtime_acl_stats_index}: begin
        acl_metadata$racl_redirect <= 'h1;
        acl_metadata$racl_nexthop <= runtime_nexthop_index;
        acl_metadata$racl_nexthop_type <= 'h0;
        acl_metadata$acl_stats_index <= runtime_acl_stats_index;
        acl_metadata$acl_copy <= runtime_acl_copy;
        fabric_metadata$reason_code <= runtime_acl_copy_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule racl_redirect_nexthop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RaclRedirectNexthopRspT {pkt: pkt, acl_metadata$racl_nexthop: acl_metadata$racl_nexthop, acl_metadata$acl_copy: acl_metadata$acl_copy, acl_metadata$acl_stats_index: acl_metadata$acl_stats_index, acl_metadata$racl_redirect: acl_metadata$racl_redirect, fabric_metadata$reason_code: fabric_metadata$reason_code, acl_metadata$racl_nexthop_type: acl_metadata$racl_nexthop_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REDIRECT_TO_CPU ======

interface RedirectToCpu;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRedirectToCpu  (RedirectToCpu);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule redirect_to_cpu_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RedirectToCpuReqT {pkt: .pkt, runtime_reason_code: .runtime_reason_code}: begin
        fabric_metadata$reason_code <= runtime_reason_code;
        fabric_metadata$dst_device <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule redirect_to_cpu_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RedirectToCpuRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, fabric_metadata$reason_code: fabric_metadata$reason_code};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REMOVE_VLAN_DOUBLE_TAGGED ======

interface RemoveVlanDoubleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRemoveVlanDoubleTagged  (RemoveVlanDoubleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule remove_vlan_double_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RemoveVlanDoubleTaggedReqT {pkt: .pkt, vlan_tag_1$etherType: .vlan_tag_1$etherType}: begin
        ethernet$etherType <= vlan_tag_1$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule remove_vlan_double_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RemoveVlanDoubleTaggedRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REMOVE_VLAN_SINGLE_TAGGED ======

interface RemoveVlanSingleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRemoveVlanSingleTagged  (RemoveVlanSingleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule remove_vlan_single_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RemoveVlanSingleTaggedReqT {pkt: .pkt, vlan_tag_0$etherType: .vlan_tag_0$etherType}: begin
        ethernet$etherType <= vlan_tag_0$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule remove_vlan_single_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RemoveVlanSingleTaggedRspT {pkt: pkt, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_IPV4_MULTICAST ======

interface RewriteIpv4Multicast;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteIpv4Multicast  (RewriteIpv4Multicast);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) ethernet$dstAddr <- mkReg(0);
  rule rewrite_ipv4_multicast_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteIpv4MulticastReqT {pkt: .pkt}: begin
        ethernet$dstAddr <= type$value;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_ipv4_multicast_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteIpv4MulticastRspT {pkt: pkt, ethernet$dstAddr: ethernet$dstAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_IPV6_MULTICAST ======

interface RewriteIpv6Multicast;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteIpv6Multicast  (RewriteIpv6Multicast);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule rewrite_ipv6_multicast_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteIpv6MulticastReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_ipv6_multicast_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteIpv6MulticastRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_SMAC ======

interface RewriteSmac;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteSmac  (RewriteSmac);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) ethernet$srcAddr <- mkReg(0);
  rule rewrite_smac_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteSmacReqT {pkt: .pkt, runtime_smac: .runtime_smac}: begin
        ethernet$srcAddr <= runtime_smac;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_smac_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteSmacRspT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_TUNNEL_DMAC ======

interface RewriteTunnelDmac;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteTunnelDmac  (RewriteTunnelDmac);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) ethernet$dstAddr <- mkReg(0);
  rule rewrite_tunnel_dmac_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteTunnelDmacReqT {pkt: .pkt, runtime_dmac: .runtime_dmac}: begin
        ethernet$dstAddr <= runtime_dmac;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_tunnel_dmac_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteTunnelDmacRspT {pkt: pkt, ethernet$dstAddr: ethernet$dstAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_TUNNEL_IPV4_DST ======

interface RewriteTunnelIpv4Dst;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteTunnelIpv4Dst  (RewriteTunnelIpv4Dst);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(32)) ipv4$dstAddr <- mkReg(0);
  rule rewrite_tunnel_ipv4_dst_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteTunnelIpv4DstReqT {pkt: .pkt, runtime_ip: .runtime_ip}: begin
        ipv4$dstAddr <= runtime_ip;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_tunnel_ipv4_dst_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteTunnelIpv4DstRspT {pkt: pkt, ipv4$dstAddr: ipv4$dstAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_TUNNEL_IPV4_SRC ======

interface RewriteTunnelIpv4Src;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteTunnelIpv4Src  (RewriteTunnelIpv4Src);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(32)) ipv4$srcAddr <- mkReg(0);
  rule rewrite_tunnel_ipv4_src_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteTunnelIpv4SrcReqT {pkt: .pkt, runtime_ip: .runtime_ip}: begin
        ipv4$srcAddr <= runtime_ip;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_tunnel_ipv4_src_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteTunnelIpv4SrcRspT {pkt: pkt, ipv4$srcAddr: ipv4$srcAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_TUNNEL_IPV6_DST ======

interface RewriteTunnelIpv6Dst;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteTunnelIpv6Dst  (RewriteTunnelIpv6Dst);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(128)) ipv6$dstAddr <- mkReg(0);
  rule rewrite_tunnel_ipv6_dst_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteTunnelIpv6DstReqT {pkt: .pkt, runtime_ip: .runtime_ip}: begin
        ipv6$dstAddr <= runtime_ip;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_tunnel_ipv6_dst_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteTunnelIpv6DstRspT {pkt: pkt, ipv6$dstAddr: ipv6$dstAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_TUNNEL_IPV6_SRC ======

interface RewriteTunnelIpv6Src;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteTunnelIpv6Src  (RewriteTunnelIpv6Src);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(128)) ipv6$srcAddr <- mkReg(0);
  rule rewrite_tunnel_ipv6_src_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteTunnelIpv6SrcReqT {pkt: .pkt, runtime_ip: .runtime_ip}: begin
        ipv6$srcAddr <= runtime_ip;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_tunnel_ipv6_src_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteTunnelIpv6SrcRspT {pkt: pkt, ipv6$srcAddr: ipv6$srcAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== REWRITE_TUNNEL_SMAC ======

interface RewriteTunnelSmac;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRewriteTunnelSmac  (RewriteTunnelSmac);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(48)) ethernet$srcAddr <- mkReg(0);
  rule rewrite_tunnel_smac_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RewriteTunnelSmacReqT {pkt: .pkt, runtime_smac: .runtime_smac}: begin
        ethernet$srcAddr <= runtime_smac;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rewrite_tunnel_smac_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RewriteTunnelSmacRspT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== RMAC_HIT ======

interface RmacHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRmacHit  (RmacHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$rmac_hit <- mkReg(0);
  rule rmac_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RmacHitReqT {pkt: .pkt}: begin
        l3_metadata$rmac_hit <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rmac_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RmacHitRspT {pkt: pkt, l3_metadata$rmac_hit: l3_metadata$rmac_hit};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== RMAC_MISS ======

interface RmacMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkRmacMiss  (RmacMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$rmac_hit <- mkReg(0);
  rule rmac_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged RmacMissReqT {pkt: .pkt}: begin
        l3_metadata$rmac_hit <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule rmac_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged RmacMissRspT {pkt: pkt, l3_metadata$rmac_hit: l3_metadata$rmac_hit};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_ACL_REDIRECT_ACTION ======

interface SetAclRedirectAction;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetAclRedirectAction  (SetAclRedirectAction);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  Reg#(Bit#(1)) nexthop_metadata$nexthop_type <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule set_acl_redirect_action_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetAclRedirectActionReqT {pkt: .pkt, acl_metadata$acl_nexthop: .acl_metadata$acl_nexthop, acl_metadata$acl_nexthop_type: .acl_metadata$acl_nexthop_type}: begin
        l3_metadata$nexthop_index <= acl_metadata$acl_nexthop;
        nexthop_metadata$nexthop_type <= acl_metadata$acl_nexthop_type;
        ingress_metadata$egress_ifindex <= 'h0;
        intrinsic_metadata$mcast_grp <= 'h0;
        fabric_metadata$dst_device <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_acl_redirect_action_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetAclRedirectActionRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, nexthop_metadata$nexthop_type: nexthop_metadata$nexthop_type, fabric_metadata$dst_device: fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_BD_FLOOD_MC_INDEX ======

interface SetBdFloodMcIndex;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetBdFloodMcIndex  (SetBdFloodMcIndex);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  rule set_bd_flood_mc_index_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetBdFloodMcIndexReqT {pkt: .pkt, runtime_mc_index: .runtime_mc_index}: begin
        intrinsic_metadata$mcast_grp <= runtime_mc_index;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_bd_flood_mc_index_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetBdFloodMcIndexRspT {pkt: pkt, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_BD_PROPERTIES ======

interface SetBdProperties;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetBdProperties  (SetBdProperties);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ingress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$outer_bd <- mkReg(0);
  Reg#(Bit#(16)) acl_metadata$bd_label <- mkReg(0);
  Reg#(Bit#(10)) l2_metadata$stp_group <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$bd_stats_idx <- mkReg(0);
  Reg#(Bit#(1)) l2_metadata$learning_enabled <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$vrf <- mkReg(0);
  Reg#(Bit#(1)) ipv4_metadata$ipv4_unicast_enabled <- mkReg(0);
  Reg#(Bit#(1)) ipv6_metadata$ipv6_unicast_enabled <- mkReg(0);
  Reg#(Bit#(2)) ipv4_metadata$ipv4_urpf_mode <- mkReg(0);
  Reg#(Bit#(2)) ipv6_metadata$ipv6_urpf_mode <- mkReg(0);
  Reg#(Bit#(10)) l3_metadata$rmac_group <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$igmp_snooping_enabled <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$mld_snooping_enabled <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$ipv4_multicast_enabled <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$ipv6_multicast_enabled <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$bd_mrpf_group <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$ipv4_mcast_key_type <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$ipv4_mcast_key <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$ipv6_mcast_key_type <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$ipv6_mcast_key <- mkReg(0);
  rule set_bd_properties_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetBdPropertiesReqT {pkt: .pkt, runtime_ipv4_multicast_enabled: .runtime_ipv4_multicast_enabled, runtime_igmp_snooping_enabled: .runtime_igmp_snooping_enabled, runtime_ipv6_mcast_key: .runtime_ipv6_mcast_key, runtime_mrpf_group: .runtime_mrpf_group, runtime_ipv4_mcast_key_type: .runtime_ipv4_mcast_key_type, runtime_mld_snooping_enabled: .runtime_mld_snooping_enabled, runtime_ipv6_multicast_enabled: .runtime_ipv6_multicast_enabled, runtime_stats_idx: .runtime_stats_idx, runtime_ipv6_urpf_mode: .runtime_ipv6_urpf_mode, runtime_ipv4_urpf_mode: .runtime_ipv4_urpf_mode, runtime_ipv4_mcast_key: .runtime_ipv4_mcast_key, runtime_bd: .runtime_bd, runtime_vrf: .runtime_vrf, runtime_learning_enabled: .runtime_learning_enabled, runtime_ipv6_unicast_enabled: .runtime_ipv6_unicast_enabled, runtime_bd_label: .runtime_bd_label, runtime_ipv6_mcast_key_type: .runtime_ipv6_mcast_key_type, runtime_rmac_group: .runtime_rmac_group, runtime_ipv4_unicast_enabled: .runtime_ipv4_unicast_enabled, runtime_stp_group: .runtime_stp_group}: begin
        ingress_metadata$bd <= runtime_bd;
        ingress_metadata$outer_bd <= runtime_bd;
        acl_metadata$bd_label <= runtime_bd_label;
        l2_metadata$stp_group <= runtime_stp_group;
        l2_metadata$bd_stats_idx <= runtime_stats_idx;
        l2_metadata$learning_enabled <= runtime_learning_enabled;
        l3_metadata$vrf <= runtime_vrf;
        ipv4_metadata$ipv4_unicast_enabled <= runtime_ipv4_unicast_enabled;
        ipv6_metadata$ipv6_unicast_enabled <= runtime_ipv6_unicast_enabled;
        ipv4_metadata$ipv4_urpf_mode <= runtime_ipv4_urpf_mode;
        ipv6_metadata$ipv6_urpf_mode <= runtime_ipv6_urpf_mode;
        l3_metadata$rmac_group <= runtime_rmac_group;
        multicast_metadata$igmp_snooping_enabled <= runtime_igmp_snooping_enabled;
        multicast_metadata$mld_snooping_enabled <= runtime_mld_snooping_enabled;
        multicast_metadata$ipv4_multicast_enabled <= runtime_ipv4_multicast_enabled;
        multicast_metadata$ipv6_multicast_enabled <= runtime_ipv6_multicast_enabled;
        multicast_metadata$bd_mrpf_group <= runtime_mrpf_group;
        multicast_metadata$ipv4_mcast_key_type <= runtime_ipv4_mcast_key_type;
        multicast_metadata$ipv4_mcast_key <= runtime_ipv4_mcast_key;
        multicast_metadata$ipv6_mcast_key_type <= runtime_ipv6_mcast_key_type;
        multicast_metadata$ipv6_mcast_key <= runtime_ipv6_mcast_key;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_bd_properties_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetBdPropertiesRspT {pkt: pkt, multicast_metadata$ipv4_mcast_key: multicast_metadata$ipv4_mcast_key, l3_metadata$rmac_group: l3_metadata$rmac_group, multicast_metadata$igmp_snooping_enabled: multicast_metadata$igmp_snooping_enabled, multicast_metadata$bd_mrpf_group: multicast_metadata$bd_mrpf_group, multicast_metadata$ipv4_multicast_enabled: multicast_metadata$ipv4_multicast_enabled, multicast_metadata$mld_snooping_enabled: multicast_metadata$mld_snooping_enabled, acl_metadata$bd_label: acl_metadata$bd_label, l2_metadata$stp_group: l2_metadata$stp_group, l3_metadata$vrf: l3_metadata$vrf, ipv6_metadata$ipv6_urpf_mode: ipv6_metadata$ipv6_urpf_mode, ipv6_metadata$ipv6_unicast_enabled: ipv6_metadata$ipv6_unicast_enabled, l2_metadata$learning_enabled: l2_metadata$learning_enabled, ingress_metadata$outer_bd: ingress_metadata$outer_bd, multicast_metadata$ipv6_mcast_key: multicast_metadata$ipv6_mcast_key, ingress_metadata$bd: ingress_metadata$bd, multicast_metadata$ipv4_mcast_key_type: multicast_metadata$ipv4_mcast_key_type, multicast_metadata$ipv6_mcast_key_type: multicast_metadata$ipv6_mcast_key_type, ipv4_metadata$ipv4_urpf_mode: ipv4_metadata$ipv4_urpf_mode, multicast_metadata$ipv6_multicast_enabled: multicast_metadata$ipv6_multicast_enabled, l2_metadata$bd_stats_idx: l2_metadata$bd_stats_idx, ipv4_metadata$ipv4_unicast_enabled: ipv4_metadata$ipv4_unicast_enabled};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_BROADCAST ======

interface SetBroadcast;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetBroadcast  (SetBroadcast);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  rule set_broadcast_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetBroadcastReqT {pkt: .pkt}: begin
        l2_metadata$lkp_pkt_type <= 'h4;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_broadcast_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetBroadcastRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$bd_stats_idx: l2_metadata$bd_stats_idx};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_CONFIG_PARAMETERS ======

interface SetConfigParameters;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetConfigParameters  (SetConfigParameters);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) intrinsic_metadata$deflect_on_drop <- mkReg(0);
  Reg#(Bit#(32)) i2e_metadata$ingress_tstamp <- mkReg(0);
  Reg#(Bit#(9)) ingress_metadata$ingress_port <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$same_if_check <- mkReg(0);
  Reg#(Bit#(9)) standard_metadata$egress_spec <- mkReg(0);
  rule set_config_parameters_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetConfigParametersReqT {pkt: .pkt, ingress_metadata$ifindex: .ingress_metadata$ifindex, intrinsic_metadata$ingress_global_tstamp: .intrinsic_metadata$ingress_global_tstamp, standard_metadata$ingress_port: .standard_metadata$ingress_port, runtime_enable_dod: .runtime_enable_dod}: begin
        intrinsic_metadata$deflect_on_drop <= runtime_enable_dod;
        i2e_metadata$ingress_tstamp <= intrinsic_metadata$ingress_global_tstamp;
        ingress_metadata$ingress_port <= standard_metadata$ingress_port;
        l2_metadata$same_if_check <= ingress_metadata$ifindex;
        standard_metadata$egress_spec <= 'h1ff;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_config_parameters_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetConfigParametersRspT {pkt: pkt, intrinsic_metadata$deflect_on_drop: intrinsic_metadata$deflect_on_drop, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp, ingress_metadata$ingress_port: ingress_metadata$ingress_port, standard_metadata$egress_spec: standard_metadata$egress_spec, l2_metadata$same_if_check: l2_metadata$same_if_check};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_CPU_REDIRECT_ACTION ======

interface SetCpuRedirectAction;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetCpuRedirectAction  (SetCpuRedirectAction);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(9)) standard_metadata$egress_spec <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule set_cpu_redirect_action_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetCpuRedirectActionReqT {pkt: .pkt}: begin
        l3_metadata$routed <= 'h0;
        intrinsic_metadata$mcast_grp <= 'h0;
        standard_metadata$egress_spec <= 'h40;
        ingress_metadata$egress_ifindex <= 'h0;
        fabric_metadata$dst_device <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_cpu_redirect_action_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetCpuRedirectActionRspT {pkt: pkt, l3_metadata$routed: l3_metadata$routed, fabric_metadata$dst_device: fabric_metadata$dst_device, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, standard_metadata$egress_spec: standard_metadata$egress_spec};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_ECMP_NEXTHOP_DETAILS ======

interface SetEcmpNexthopDetails;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetEcmpNexthopDetails  (SetEcmpNexthopDetails);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  rule set_ecmp_nexthop_details_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetEcmpNexthopDetailsReqT {pkt: .pkt, runtime_bd: .runtime_bd, runtime_nhop_index: .runtime_nhop_index, runtime_ifindex: .runtime_ifindex, runtime_tunnel: .runtime_tunnel}: begin
        ingress_metadata$egress_ifindex <= runtime_ifindex;
        l3_metadata$nexthop_index <= runtime_nhop_index;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_ecmp_nexthop_details_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetEcmpNexthopDetailsRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_ECMP_NEXTHOP_DETAILS_FOR_POST_ROUTED_FLOOD ======

interface SetEcmpNexthopDetailsForPostRoutedFlood;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetEcmpNexthopDetailsForPostRoutedFlood  (SetEcmpNexthopDetailsForPostRoutedFlood);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule set_ecmp_nexthop_details_for_post_routed_flood_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetEcmpNexthopDetailsForPostRoutedFloodReqT {pkt: .pkt, runtime_uuc_mc_index: .runtime_uuc_mc_index, runtime_nhop_index: .runtime_nhop_index, runtime_bd: .runtime_bd}: begin
        intrinsic_metadata$mcast_grp <= runtime_uuc_mc_index;
        l3_metadata$nexthop_index <= runtime_nhop_index;
        ingress_metadata$egress_ifindex <= 'h0;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_ecmp_nexthop_details_for_post_routed_flood_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetEcmpNexthopDetailsForPostRoutedFloodRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, fabric_metadata$dst_device: fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_EGRESS_BD_PROPERTIES ======

interface SetEgressBdProperties;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetEgressBdProperties  (SetEgressBdProperties);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(9)) egress_metadata$smac_idx <- mkReg(0);
  rule set_egress_bd_properties_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetEgressBdPropertiesReqT {pkt: .pkt, runtime_smac_idx: .runtime_smac_idx}: begin
        egress_metadata$smac_idx <= runtime_smac_idx;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_egress_bd_properties_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetEgressBdPropertiesRspT {pkt: pkt, egress_metadata$smac_idx: egress_metadata$smac_idx};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_EGRESS_FILTER_DROP ======

interface SetEgressFilterDrop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetEgressFilterDrop  (SetEgressFilterDrop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule set_egress_filter_drop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetEgressFilterDropReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_egress_filter_drop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetEgressFilterDropRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_EGRESS_PACKET_VLAN_DOUBLE_TAGGED ======

interface SetEgressPacketVlanDoubleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetEgressPacketVlanDoubleTagged  (SetEgressPacketVlanDoubleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) vlan_tag_1$etherType <- mkReg(0);
  Reg#(Bit#(12)) vlan_tag_1$vid <- mkReg(0);
  Reg#(Bit#(16)) vlan_tag_0$etherType <- mkReg(0);
  Reg#(Bit#(12)) vlan_tag_0$vid <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule set_egress_packet_vlan_double_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetEgressPacketVlanDoubleTaggedReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType, runtime_c_tag: .runtime_c_tag, runtime_s_tag: .runtime_s_tag}: begin
        vlan_tag_1$etherType <= ethernet$etherType;
        vlan_tag_1$vid <= runtime_c_tag;
        vlan_tag_0$etherType <= 'h8100;
        vlan_tag_0$vid <= runtime_s_tag;
        ethernet$etherType <= 'h9100;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_egress_packet_vlan_double_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetEgressPacketVlanDoubleTaggedRspT {pkt: pkt, vlan_tag_1$vid: vlan_tag_1$vid, vlan_tag_0$vid: vlan_tag_0$vid, vlan_tag_0$etherType: vlan_tag_0$etherType, vlan_tag_1$etherType: vlan_tag_1$etherType, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_EGRESS_PACKET_VLAN_TAGGED ======

interface SetEgressPacketVlanTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetEgressPacketVlanTagged  (SetEgressPacketVlanTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) vlan_tag_0$etherType <- mkReg(0);
  Reg#(Bit#(12)) vlan_tag_0$vid <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule set_egress_packet_vlan_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetEgressPacketVlanTaggedReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType, runtime_vlan_id: .runtime_vlan_id}: begin
        vlan_tag_0$etherType <= ethernet$etherType;
        vlan_tag_0$vid <= runtime_vlan_id;
        ethernet$etherType <= 'h8100;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_egress_packet_vlan_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetEgressPacketVlanTaggedRspT {pkt: pkt, vlan_tag_0$vid: vlan_tag_0$vid, vlan_tag_0$etherType: vlan_tag_0$etherType, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_EGRESS_PACKET_VLAN_UNTAGGED ======

interface SetEgressPacketVlanUntagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetEgressPacketVlanUntagged  (SetEgressPacketVlanUntagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule set_egress_packet_vlan_untagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetEgressPacketVlanUntaggedReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_egress_packet_vlan_untagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetEgressPacketVlanUntaggedRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_EGRESS_TUNNEL_VNI ======

interface SetEgressTunnelVni;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetEgressTunnelVni  (SetEgressTunnelVni);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(24)) tunnel_metadata$vnid <- mkReg(0);
  rule set_egress_tunnel_vni_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetEgressTunnelVniReqT {pkt: .pkt, runtime_vnid: .runtime_vnid}: begin
        tunnel_metadata$vnid <= runtime_vnid;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_egress_tunnel_vni_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetEgressTunnelVniRspT {pkt: pkt, tunnel_metadata$vnid: tunnel_metadata$vnid};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_FABRIC_LAG_PORT ======

interface SetFabricLagPort;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetFabricLagPort  (SetFabricLagPort);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(9)) standard_metadata$egress_spec <- mkReg(0);
  rule set_fabric_lag_port_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetFabricLagPortReqT {pkt: .pkt, runtime_port: .runtime_port}: begin
        standard_metadata$egress_spec <= runtime_port;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_fabric_lag_port_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetFabricLagPortRspT {pkt: pkt, standard_metadata$egress_spec: standard_metadata$egress_spec};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_FABRIC_MULTICAST ======

interface SetFabricMulticast;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetFabricMulticast  (SetFabricMulticast);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) multicast_metadata$mcast_grp <- mkReg(0);
  rule set_fabric_multicast_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetFabricMulticastReqT {pkt: .pkt, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        multicast_metadata$mcast_grp <= intrinsic_metadata$mcast_grp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_fabric_multicast_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetFabricMulticastRspT {pkt: pkt, multicast_metadata$mcast_grp: multicast_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_FIB_REDIRECT_ACTION ======

interface SetFibRedirectAction;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetFibRedirectAction  (SetFibRedirectAction);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  Reg#(Bit#(1)) nexthop_metadata$nexthop_type <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule set_fib_redirect_action_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetFibRedirectActionReqT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        l3_metadata$nexthop_index <= l3_metadata$fib_nexthop;
        nexthop_metadata$nexthop_type <= l3_metadata$fib_nexthop_type;
        l3_metadata$routed <= 'h1;
        intrinsic_metadata$mcast_grp <= 'h0;
        fabric_metadata$reason_code <= 'h217;
        fabric_metadata$dst_device <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_fib_redirect_action_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetFibRedirectActionRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, nexthop_metadata$nexthop_type: nexthop_metadata$nexthop_type, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, l3_metadata$routed: l3_metadata$routed, fabric_metadata$dst_device: fabric_metadata$dst_device, fabric_metadata$reason_code: fabric_metadata$reason_code};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_IFINDEX ======

interface SetIfindex;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetIfindex  (SetIfindex);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ingress_metadata$ifindex <- mkReg(0);
  Reg#(Bit#(2)) ingress_metadata$port_type <- mkReg(0);
  rule set_ifindex_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetIfindexReqT {pkt: .pkt, runtime_port_type: .runtime_port_type, runtime_ifindex: .runtime_ifindex}: begin
        ingress_metadata$ifindex <= runtime_ifindex;
        ingress_metadata$port_type <= runtime_port_type;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_ifindex_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetIfindexRspT {pkt: pkt, ingress_metadata$port_type: ingress_metadata$port_type, ingress_metadata$ifindex: ingress_metadata$ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_INGRESS_IFINDEX_PROPERTIES ======

interface SetIngressIfindexProperties;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetIngressIfindexProperties  (SetIngressIfindexProperties);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule set_ingress_ifindex_properties_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetIngressIfindexPropertiesReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_ingress_ifindex_properties_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetIngressIfindexPropertiesRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_INGRESS_PORT_PROPERTIES ======

interface SetIngressPortProperties;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetIngressPortProperties  (SetIngressPortProperties);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) acl_metadata$if_label <- mkReg(0);
  rule set_ingress_port_properties_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetIngressPortPropertiesReqT {pkt: .pkt, runtime_if_label: .runtime_if_label}: begin
        acl_metadata$if_label <= runtime_if_label;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_ingress_port_properties_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetIngressPortPropertiesRspT {pkt: pkt, acl_metadata$if_label: acl_metadata$if_label};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_L2_REDIRECT_ACTION ======

interface SetL2RedirectAction;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetL2RedirectAction  (SetL2RedirectAction);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  Reg#(Bit#(1)) nexthop_metadata$nexthop_type <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule set_l2_redirect_action_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetL2RedirectActionReqT {pkt: .pkt, l2_metadata$l2_nexthop: .l2_metadata$l2_nexthop, l2_metadata$l2_nexthop_type: .l2_metadata$l2_nexthop_type}: begin
        l3_metadata$nexthop_index <= l2_metadata$l2_nexthop;
        nexthop_metadata$nexthop_type <= l2_metadata$l2_nexthop_type;
        ingress_metadata$egress_ifindex <= 'h0;
        intrinsic_metadata$mcast_grp <= 'h0;
        fabric_metadata$dst_device <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_l2_redirect_action_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetL2RedirectActionRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, nexthop_metadata$nexthop_type: nexthop_metadata$nexthop_type, fabric_metadata$dst_device: fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_L2_REWRITE ======

interface SetL2Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetL2Rewrite  (SetL2Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$outer_bd <- mkReg(0);
  rule set_l2_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetL2RewriteReqT {pkt: .pkt, ingress_metadata$bd: .ingress_metadata$bd}: begin
        egress_metadata$routed <= 'h0;
        egress_metadata$bd <= ingress_metadata$bd;
        egress_metadata$outer_bd <= ingress_metadata$bd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_l2_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetL2RewriteRspT {pkt: pkt, egress_metadata$outer_bd: egress_metadata$outer_bd, egress_metadata$bd: egress_metadata$bd, egress_metadata$routed: egress_metadata$routed};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_L2_REWRITE_WITH_TUNNEL ======

interface SetL2RewriteWithTunnel;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetL2RewriteWithTunnel  (SetL2RewriteWithTunnel);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$outer_bd <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  rule set_l2_rewrite_with_tunnel_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetL2RewriteWithTunnelReqT {pkt: .pkt, ingress_metadata$bd: .ingress_metadata$bd, runtime_tunnel_index: .runtime_tunnel_index, runtime_tunnel_type: .runtime_tunnel_type}: begin
        egress_metadata$routed <= 'h0;
        egress_metadata$bd <= ingress_metadata$bd;
        egress_metadata$outer_bd <= ingress_metadata$bd;
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        tunnel_metadata$egress_tunnel_type <= runtime_tunnel_type;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_l2_rewrite_with_tunnel_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetL2RewriteWithTunnelRspT {pkt: pkt, egress_metadata$outer_bd: egress_metadata$outer_bd, egress_metadata$bd: egress_metadata$bd, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index, egress_metadata$routed: egress_metadata$routed, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_L3_REWRITE ======

interface SetL3Rewrite;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetL3Rewrite  (SetL3Rewrite);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(48)) egress_metadata$mac_da <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$outer_bd <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$mtu_index <- mkReg(0);
  rule set_l3_rewrite_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetL3RewriteReqT {pkt: .pkt, runtime_dmac: .runtime_dmac, runtime_bd: .runtime_bd, runtime_mtu_index: .runtime_mtu_index}: begin
        egress_metadata$routed <= 'h1;
        egress_metadata$mac_da <= runtime_dmac;
        egress_metadata$bd <= runtime_bd;
        egress_metadata$outer_bd <= runtime_bd;
        l3_metadata$mtu_index <= runtime_mtu_index;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_l3_rewrite_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetL3RewriteRspT {pkt: pkt, egress_metadata$outer_bd: egress_metadata$outer_bd, egress_metadata$bd: egress_metadata$bd, egress_metadata$mac_da: egress_metadata$mac_da, egress_metadata$routed: egress_metadata$routed, l3_metadata$mtu_index: l3_metadata$mtu_index};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_L3_REWRITE_WITH_TUNNEL ======

interface SetL3RewriteWithTunnel;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetL3RewriteWithTunnel  (SetL3RewriteWithTunnel);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(48)) egress_metadata$mac_da <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$outer_bd <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  rule set_l3_rewrite_with_tunnel_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetL3RewriteWithTunnelReqT {pkt: .pkt, runtime_dmac: .runtime_dmac, runtime_tunnel_index: .runtime_tunnel_index, runtime_bd: .runtime_bd, runtime_tunnel_type: .runtime_tunnel_type}: begin
        egress_metadata$routed <= 'h1;
        egress_metadata$mac_da <= runtime_dmac;
        egress_metadata$bd <= runtime_bd;
        egress_metadata$outer_bd <= runtime_bd;
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        tunnel_metadata$egress_tunnel_type <= runtime_tunnel_type;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_l3_rewrite_with_tunnel_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetL3RewriteWithTunnelRspT {pkt: pkt, egress_metadata$outer_bd: egress_metadata$outer_bd, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index, egress_metadata$mac_da: egress_metadata$mac_da, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type, egress_metadata$bd: egress_metadata$bd, egress_metadata$routed: egress_metadata$routed};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_LAG_MISS ======

interface SetLagMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetLagMiss  (SetLagMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule set_lag_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetLagMissReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_lag_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetLagMissRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_LAG_PORT ======

interface SetLagPort;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetLagPort  (SetLagPort);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(9)) standard_metadata$egress_spec <- mkReg(0);
  rule set_lag_port_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetLagPortReqT {pkt: .pkt, runtime_port: .runtime_port}: begin
        standard_metadata$egress_spec <= runtime_port;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_lag_port_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetLagPortRspT {pkt: pkt, standard_metadata$egress_spec: standard_metadata$egress_spec};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_LAG_REMOTE_PORT ======

interface SetLagRemotePort;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetLagRemotePort  (SetLagRemotePort);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$dst_port <- mkReg(0);
  rule set_lag_remote_port_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetLagRemotePortReqT {pkt: .pkt, runtime_device: .runtime_device, runtime_port: .runtime_port}: begin
        fabric_metadata$dst_device <= runtime_device;
        fabric_metadata$dst_port <= runtime_port;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_lag_remote_port_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetLagRemotePortRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, fabric_metadata$dst_port: fabric_metadata$dst_port};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MALFORMED_OUTER_IPV4_PACKET ======

interface SetMalformedOuterIpv4Packet;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMalformedOuterIpv4Packet  (SetMalformedOuterIpv4Packet);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) ingress_metadata$drop_flag <- mkReg(0);
  Reg#(Bit#(8)) ingress_metadata$drop_reason <- mkReg(0);
  rule set_malformed_outer_ipv4_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMalformedOuterIpv4PacketReqT {pkt: .pkt, runtime_drop_reason: .runtime_drop_reason}: begin
        ingress_metadata$drop_flag <= 'h1;
        ingress_metadata$drop_reason <= runtime_drop_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_malformed_outer_ipv4_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMalformedOuterIpv4PacketRspT {pkt: pkt, ingress_metadata$drop_reason: ingress_metadata$drop_reason, ingress_metadata$drop_flag: ingress_metadata$drop_flag};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MALFORMED_OUTER_IPV6_PACKET ======

interface SetMalformedOuterIpv6Packet;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMalformedOuterIpv6Packet  (SetMalformedOuterIpv6Packet);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) ingress_metadata$drop_flag <- mkReg(0);
  Reg#(Bit#(8)) ingress_metadata$drop_reason <- mkReg(0);
  rule set_malformed_outer_ipv6_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMalformedOuterIpv6PacketReqT {pkt: .pkt, runtime_drop_reason: .runtime_drop_reason}: begin
        ingress_metadata$drop_flag <= 'h1;
        ingress_metadata$drop_reason <= runtime_drop_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_malformed_outer_ipv6_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMalformedOuterIpv6PacketRspT {pkt: pkt, ingress_metadata$drop_reason: ingress_metadata$drop_reason, ingress_metadata$drop_flag: ingress_metadata$drop_flag};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MALFORMED_PACKET ======

interface SetMalformedPacket;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMalformedPacket  (SetMalformedPacket);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) ingress_metadata$drop_flag <- mkReg(0);
  Reg#(Bit#(8)) ingress_metadata$drop_reason <- mkReg(0);
  rule set_malformed_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMalformedPacketReqT {pkt: .pkt, runtime_drop_reason: .runtime_drop_reason}: begin
        ingress_metadata$drop_flag <= 'h1;
        ingress_metadata$drop_reason <= runtime_drop_reason;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_malformed_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMalformedPacketRspT {pkt: pkt, ingress_metadata$drop_reason: ingress_metadata$drop_reason, ingress_metadata$drop_flag: ingress_metadata$drop_flag};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MIRROR_BD ======

interface SetMirrorBd;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMirrorBd  (SetMirrorBd);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  rule set_mirror_bd_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMirrorBdReqT {pkt: .pkt, runtime_bd: .runtime_bd}: begin
        egress_metadata$bd <= runtime_bd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mirror_bd_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMirrorBdRspT {pkt: pkt, egress_metadata$bd: egress_metadata$bd};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MIRROR_NHOP ======

interface SetMirrorNhop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMirrorNhop  (SetMirrorNhop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  rule set_mirror_nhop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMirrorNhopReqT {pkt: .pkt, runtime_nhop_idx: .runtime_nhop_idx}: begin
        l3_metadata$nexthop_index <= runtime_nhop_idx;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mirror_nhop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMirrorNhopRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MPLS_PUSH_REWRITE_L2 ======

interface SetMplsPushRewriteL2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMplsPushRewriteL2  (SetMplsPushRewriteL2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  Reg#(Bit#(4)) tunnel_metadata$egress_header_count <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  rule set_mpls_push_rewrite_l2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMplsPushRewriteL2ReqT {pkt: .pkt, l3_metadata$routed: .l3_metadata$routed, ingress_metadata$bd: .ingress_metadata$bd, runtime_tunnel_index: .runtime_tunnel_index, runtime_header_count: .runtime_header_count}: begin
        egress_metadata$routed <= l3_metadata$routed;
        egress_metadata$bd <= ingress_metadata$bd;
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        tunnel_metadata$egress_header_count <= runtime_header_count;
        tunnel_metadata$egress_tunnel_type <= 'hd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mpls_push_rewrite_l2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMplsPushRewriteL2RspT {pkt: pkt, egress_metadata$bd: egress_metadata$bd, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index, tunnel_metadata$egress_header_count: tunnel_metadata$egress_header_count, egress_metadata$routed: egress_metadata$routed, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MPLS_PUSH_REWRITE_L3 ======

interface SetMplsPushRewriteL3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMplsPushRewriteL3  (SetMplsPushRewriteL3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(48)) egress_metadata$mac_da <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  Reg#(Bit#(4)) tunnel_metadata$egress_header_count <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  rule set_mpls_push_rewrite_l3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMplsPushRewriteL3ReqT {pkt: .pkt, l3_metadata$routed: .l3_metadata$routed, runtime_dmac: .runtime_dmac, runtime_tunnel_index: .runtime_tunnel_index, runtime_bd: .runtime_bd, runtime_header_count: .runtime_header_count}: begin
        egress_metadata$routed <= l3_metadata$routed;
        egress_metadata$bd <= runtime_bd;
        egress_metadata$mac_da <= runtime_dmac;
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        tunnel_metadata$egress_header_count <= runtime_header_count;
        tunnel_metadata$egress_tunnel_type <= 'he;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mpls_push_rewrite_l3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMplsPushRewriteL3RspT {pkt: pkt, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index, egress_metadata$routed: egress_metadata$routed, egress_metadata$mac_da: egress_metadata$mac_da, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type, egress_metadata$bd: egress_metadata$bd, tunnel_metadata$egress_header_count: tunnel_metadata$egress_header_count};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MPLS_REWRITE_PUSH1 ======

interface SetMplsRewritePush1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMplsRewritePush1  (SetMplsRewritePush1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(20)) mpls0$label <- mkReg(0);
  Reg#(Bit#(3)) mpls0$exp <- mkReg(0);
  Reg#(Bit#(1)) mpls0$bos <- mkReg(0);
  Reg#(Bit#(8)) mpls0$ttl <- mkReg(0);
  Reg#(Bit#(9)) tunnel_metadata$tunnel_smac_index <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_dmac_index <- mkReg(0);
  rule set_mpls_rewrite_push1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMplsRewritePush1ReqT {pkt: .pkt, runtime_ttl1: .runtime_ttl1, runtime_exp1: .runtime_exp1, runtime_label1: .runtime_label1, runtime_dmac_idx: .runtime_dmac_idx, runtime_smac_idx: .runtime_smac_idx}: begin
        mpls0$label <= runtime_label1;
        mpls0$exp <= runtime_exp1;
        mpls0$bos <= 'h1;
        mpls0$ttl <= runtime_ttl1;
        tunnel_metadata$tunnel_smac_index <= runtime_smac_idx;
        tunnel_metadata$tunnel_dmac_index <= runtime_dmac_idx;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mpls_rewrite_push1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMplsRewritePush1RspT {pkt: pkt, tunnel_metadata$tunnel_smac_index: tunnel_metadata$tunnel_smac_index, mpls0$exp: mpls0$exp, mpls0$ttl: mpls0$ttl, mpls0$bos: mpls0$bos, tunnel_metadata$tunnel_dmac_index: tunnel_metadata$tunnel_dmac_index, mpls0$label: mpls0$label};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MPLS_REWRITE_PUSH2 ======

interface SetMplsRewritePush2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMplsRewritePush2  (SetMplsRewritePush2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(20)) mpls0$label <- mkReg(0);
  Reg#(Bit#(3)) mpls0$exp <- mkReg(0);
  Reg#(Bit#(8)) mpls0$ttl <- mkReg(0);
  Reg#(Bit#(1)) mpls0$bos <- mkReg(0);
  Reg#(Bit#(20)) mpls1$label <- mkReg(0);
  Reg#(Bit#(3)) mpls1$exp <- mkReg(0);
  Reg#(Bit#(8)) mpls1$ttl <- mkReg(0);
  Reg#(Bit#(1)) mpls1$bos <- mkReg(0);
  Reg#(Bit#(9)) tunnel_metadata$tunnel_smac_index <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_dmac_index <- mkReg(0);
  rule set_mpls_rewrite_push2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMplsRewritePush2ReqT {pkt: .pkt, runtime_exp1: .runtime_exp1, runtime_ttl2: .runtime_ttl2, runtime_smac_idx: .runtime_smac_idx, runtime_ttl1: .runtime_ttl1, runtime_label2: .runtime_label2, runtime_exp2: .runtime_exp2, runtime_label1: .runtime_label1, runtime_dmac_idx: .runtime_dmac_idx}: begin
        mpls0$label <= runtime_label1;
        mpls0$exp <= runtime_exp1;
        mpls0$ttl <= runtime_ttl1;
        mpls0$bos <= 'h0;
        mpls1$label <= runtime_label2;
        mpls1$exp <= runtime_exp2;
        mpls1$ttl <= runtime_ttl2;
        mpls1$bos <= 'h1;
        tunnel_metadata$tunnel_smac_index <= runtime_smac_idx;
        tunnel_metadata$tunnel_dmac_index <= runtime_dmac_idx;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mpls_rewrite_push2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMplsRewritePush2RspT {pkt: pkt, mpls1$ttl: mpls1$ttl, tunnel_metadata$tunnel_smac_index: tunnel_metadata$tunnel_smac_index, mpls1$exp: mpls1$exp, mpls0$exp: mpls0$exp, mpls0$ttl: mpls0$ttl, mpls1$label: mpls1$label, mpls0$bos: mpls0$bos, mpls1$bos: mpls1$bos, tunnel_metadata$tunnel_dmac_index: tunnel_metadata$tunnel_dmac_index, mpls0$label: mpls0$label};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MPLS_REWRITE_PUSH3 ======

interface SetMplsRewritePush3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMplsRewritePush3  (SetMplsRewritePush3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(20)) mpls0$label <- mkReg(0);
  Reg#(Bit#(3)) mpls0$exp <- mkReg(0);
  Reg#(Bit#(8)) mpls0$ttl <- mkReg(0);
  Reg#(Bit#(1)) mpls0$bos <- mkReg(0);
  Reg#(Bit#(20)) mpls1$label <- mkReg(0);
  Reg#(Bit#(3)) mpls1$exp <- mkReg(0);
  Reg#(Bit#(8)) mpls1$ttl <- mkReg(0);
  Reg#(Bit#(1)) mpls1$bos <- mkReg(0);
  Reg#(Bit#(20)) mpls2$label <- mkReg(0);
  Reg#(Bit#(3)) mpls2$exp <- mkReg(0);
  Reg#(Bit#(8)) mpls2$ttl <- mkReg(0);
  Reg#(Bit#(1)) mpls2$bos <- mkReg(0);
  Reg#(Bit#(9)) tunnel_metadata$tunnel_smac_index <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_dmac_index <- mkReg(0);
  rule set_mpls_rewrite_push3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMplsRewritePush3ReqT {pkt: .pkt, runtime_exp3: .runtime_exp3, runtime_exp1: .runtime_exp1, runtime_ttl2: .runtime_ttl2, runtime_label3: .runtime_label3, runtime_ttl1: .runtime_ttl1, runtime_label2: .runtime_label2, runtime_exp2: .runtime_exp2, runtime_label1: .runtime_label1, runtime_smac_idx: .runtime_smac_idx, runtime_ttl3: .runtime_ttl3, runtime_dmac_idx: .runtime_dmac_idx}: begin
        mpls0$label <= runtime_label1;
        mpls0$exp <= runtime_exp1;
        mpls0$ttl <= runtime_ttl1;
        mpls0$bos <= 'h0;
        mpls1$label <= runtime_label2;
        mpls1$exp <= runtime_exp2;
        mpls1$ttl <= runtime_ttl2;
        mpls1$bos <= 'h0;
        mpls2$label <= runtime_label3;
        mpls2$exp <= runtime_exp3;
        mpls2$ttl <= runtime_ttl3;
        mpls2$bos <= 'h1;
        tunnel_metadata$tunnel_smac_index <= runtime_smac_idx;
        tunnel_metadata$tunnel_dmac_index <= runtime_dmac_idx;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mpls_rewrite_push3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMplsRewritePush3RspT {pkt: pkt, mpls1$ttl: mpls1$ttl, mpls1$exp: mpls1$exp, mpls2$bos: mpls2$bos, tunnel_metadata$tunnel_smac_index: tunnel_metadata$tunnel_smac_index, mpls1$label: mpls1$label, mpls0$bos: mpls0$bos, mpls2$exp: mpls2$exp, mpls2$ttl: mpls2$ttl, mpls0$exp: mpls0$exp, tunnel_metadata$tunnel_dmac_index: tunnel_metadata$tunnel_dmac_index, mpls0$ttl: mpls0$ttl, mpls2$label: mpls2$label, mpls1$bos: mpls1$bos, mpls0$label: mpls0$label};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MPLS_SWAP_PUSH_REWRITE_L2 ======

interface SetMplsSwapPushRewriteL2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMplsSwapPushRewriteL2  (SetMplsSwapPushRewriteL2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(20)) mpls0$label <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  Reg#(Bit#(4)) tunnel_metadata$egress_header_count <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  rule set_mpls_swap_push_rewrite_l2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMplsSwapPushRewriteL2ReqT {pkt: .pkt, l3_metadata$routed: .l3_metadata$routed, ingress_metadata$bd: .ingress_metadata$bd, runtime_tunnel_index: .runtime_tunnel_index, runtime_label: .runtime_label, runtime_header_count: .runtime_header_count}: begin
        egress_metadata$routed <= l3_metadata$routed;
        egress_metadata$bd <= ingress_metadata$bd;
        mpls0$label <= runtime_label;
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        tunnel_metadata$egress_header_count <= runtime_header_count;
        tunnel_metadata$egress_tunnel_type <= 'hd;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mpls_swap_push_rewrite_l2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMplsSwapPushRewriteL2RspT {pkt: pkt, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index, egress_metadata$routed: egress_metadata$routed, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type, egress_metadata$bd: egress_metadata$bd, tunnel_metadata$egress_header_count: tunnel_metadata$egress_header_count, mpls0$label: mpls0$label};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MPLS_SWAP_PUSH_REWRITE_L3 ======

interface SetMplsSwapPushRewriteL3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMplsSwapPushRewriteL3  (SetMplsSwapPushRewriteL3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) egress_metadata$bd <- mkReg(0);
  Reg#(Bit#(20)) mpls0$label <- mkReg(0);
  Reg#(Bit#(48)) egress_metadata$mac_da <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_index <- mkReg(0);
  Reg#(Bit#(4)) tunnel_metadata$egress_header_count <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$egress_tunnel_type <- mkReg(0);
  rule set_mpls_swap_push_rewrite_l3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMplsSwapPushRewriteL3ReqT {pkt: .pkt, l3_metadata$routed: .l3_metadata$routed, runtime_dmac: .runtime_dmac, runtime_tunnel_index: .runtime_tunnel_index, runtime_label: .runtime_label, runtime_bd: .runtime_bd, runtime_header_count: .runtime_header_count}: begin
        egress_metadata$routed <= l3_metadata$routed;
        egress_metadata$bd <= runtime_bd;
        mpls0$label <= runtime_label;
        egress_metadata$mac_da <= runtime_dmac;
        tunnel_metadata$tunnel_index <= runtime_tunnel_index;
        tunnel_metadata$egress_header_count <= runtime_header_count;
        tunnel_metadata$egress_tunnel_type <= 'he;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_mpls_swap_push_rewrite_l3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMplsSwapPushRewriteL3RspT {pkt: pkt, tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index, tunnel_metadata$egress_header_count: tunnel_metadata$egress_header_count, egress_metadata$mac_da: egress_metadata$mac_da, tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type, egress_metadata$bd: egress_metadata$bd, egress_metadata$routed: egress_metadata$routed, mpls0$label: mpls0$label};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MULTICAST ======

interface SetMulticast;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMulticast  (SetMulticast);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  rule set_multicast_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMulticastReqT {pkt: .pkt}: begin
        l2_metadata$lkp_pkt_type <= 'h2;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_multicast_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMulticastRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$bd_stats_idx: l2_metadata$bd_stats_idx};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MULTICAST_AND_IPV6_SRC_IS_LINK_LOCAL ======

interface SetMulticastAndIpv6SrcIsLinkLocal;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMulticastAndIpv6SrcIsLinkLocal  (SetMulticastAndIpv6SrcIsLinkLocal);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(1)) ipv6_metadata$ipv6_src_is_link_local <- mkReg(0);
  rule set_multicast_and_ipv6_src_is_link_local_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMulticastAndIpv6SrcIsLinkLocalReqT {pkt: .pkt}: begin
        l2_metadata$lkp_pkt_type <= 'h2;
        ipv6_metadata$ipv6_src_is_link_local <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_multicast_and_ipv6_src_is_link_local_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMulticastAndIpv6SrcIsLinkLocalRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, ipv6_metadata$ipv6_src_is_link_local: ipv6_metadata$ipv6_src_is_link_local, l2_metadata$bd_stats_idx: l2_metadata$bd_stats_idx};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MULTICAST_BRIDGE_ACTION ======

interface SetMulticastBridgeAction;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMulticastBridgeAction  (SetMulticastBridgeAction);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  rule set_multicast_bridge_action_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMulticastBridgeActionReqT {pkt: .pkt, multicast_metadata$multicast_bridge_mc_index: .multicast_metadata$multicast_bridge_mc_index}: begin
        fabric_metadata$dst_device <= 'h7f;
        ingress_metadata$egress_ifindex <= 'h0;
        intrinsic_metadata$mcast_grp <= multicast_metadata$multicast_bridge_mc_index;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_multicast_bridge_action_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMulticastBridgeActionRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MULTICAST_DROP ======

interface SetMulticastDrop;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMulticastDrop  (SetMulticastDrop);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) ingress_metadata$drop_flag <- mkReg(0);
  Reg#(Bit#(8)) ingress_metadata$drop_reason <- mkReg(0);
  rule set_multicast_drop_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMulticastDropReqT {pkt: .pkt}: begin
        ingress_metadata$drop_flag <= 'h1;
        ingress_metadata$drop_reason <= 'h2c;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_multicast_drop_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMulticastDropRspT {pkt: pkt, ingress_metadata$drop_reason: ingress_metadata$drop_reason, ingress_metadata$drop_flag: ingress_metadata$drop_flag};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MULTICAST_FLOOD ======

interface SetMulticastFlood;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMulticastFlood  (SetMulticastFlood);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  rule set_multicast_flood_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMulticastFloodReqT {pkt: .pkt}: begin
        fabric_metadata$dst_device <= 'h7f;
        ingress_metadata$egress_ifindex <= 'hffff;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_multicast_flood_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMulticastFloodRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_MULTICAST_ROUTE_ACTION ======

interface SetMulticastRouteAction;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetMulticastRouteAction  (SetMulticastRouteAction);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$same_bd_check <- mkReg(0);
  rule set_multicast_route_action_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetMulticastRouteActionReqT {pkt: .pkt, multicast_metadata$multicast_route_mc_index: .multicast_metadata$multicast_route_mc_index}: begin
        fabric_metadata$dst_device <= 'h7f;
        ingress_metadata$egress_ifindex <= 'h0;
        intrinsic_metadata$mcast_grp <= multicast_metadata$multicast_route_mc_index;
        l3_metadata$routed <= 'h1;
        l3_metadata$same_bd_check <= 'hffff;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_multicast_route_action_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetMulticastRouteActionRspT {pkt: pkt, l3_metadata$routed: l3_metadata$routed, fabric_metadata$dst_device: fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, l3_metadata$same_bd_check: l3_metadata$same_bd_check, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_NEXTHOP_DETAILS ======

interface SetNexthopDetails;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetNexthopDetails  (SetNexthopDetails);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  rule set_nexthop_details_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetNexthopDetailsReqT {pkt: .pkt, runtime_bd: .runtime_bd, runtime_tunnel: .runtime_tunnel, runtime_ifindex: .runtime_ifindex}: begin
        ingress_metadata$egress_ifindex <= runtime_ifindex;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_nexthop_details_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetNexthopDetailsRspT {pkt: pkt, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_NEXTHOP_DETAILS_FOR_POST_ROUTED_FLOOD ======

interface SetNexthopDetailsForPostRoutedFlood;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetNexthopDetailsForPostRoutedFlood  (SetNexthopDetailsForPostRoutedFlood);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule set_nexthop_details_for_post_routed_flood_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetNexthopDetailsForPostRoutedFloodReqT {pkt: .pkt, runtime_uuc_mc_index: .runtime_uuc_mc_index, runtime_bd: .runtime_bd}: begin
        intrinsic_metadata$mcast_grp <= runtime_uuc_mc_index;
        ingress_metadata$egress_ifindex <= 'h0;
        fabric_metadata$dst_device <= 'h7f;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_nexthop_details_for_post_routed_flood_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetNexthopDetailsForPostRoutedFloodRspT {pkt: pkt, fabric_metadata$dst_device: fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_RACL_REDIRECT_ACTION ======

interface SetRaclRedirectAction;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetRaclRedirectAction  (SetRaclRedirectAction);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  Reg#(Bit#(1)) nexthop_metadata$nexthop_type <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$routed <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  rule set_racl_redirect_action_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetRaclRedirectActionReqT {pkt: .pkt, acl_metadata$racl_nexthop: .acl_metadata$racl_nexthop, acl_metadata$racl_nexthop_type: .acl_metadata$racl_nexthop_type}: begin
        l3_metadata$nexthop_index <= acl_metadata$racl_nexthop;
        nexthop_metadata$nexthop_type <= acl_metadata$racl_nexthop_type;
        l3_metadata$routed <= 'h1;
        ingress_metadata$egress_ifindex <= 'h0;
        intrinsic_metadata$mcast_grp <= 'h0;
        fabric_metadata$dst_device <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_racl_redirect_action_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetRaclRedirectActionRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, nexthop_metadata$nexthop_type: nexthop_metadata$nexthop_type, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex, l3_metadata$routed: l3_metadata$routed, fabric_metadata$dst_device: fabric_metadata$dst_device};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_REPLICA_COPY_BRIDGED ======

interface SetReplicaCopyBridged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetReplicaCopyBridged  (SetReplicaCopyBridged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) egress_metadata$routed <- mkReg(0);
  rule set_replica_copy_bridged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetReplicaCopyBridgedReqT {pkt: .pkt}: begin
        egress_metadata$routed <= 'h0;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_replica_copy_bridged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetReplicaCopyBridgedRspT {pkt: pkt, egress_metadata$routed: egress_metadata$routed};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_STORM_CONTROL_METER ======

interface SetStormControlMeter;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetStormControlMeter  (SetStormControlMeter);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) meter_metadata$meter_index <- mkReg(0);
  rule set_storm_control_meter_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetStormControlMeterReqT {pkt: .pkt, runtime_meter_idx: .runtime_meter_idx}: begin
        meter_metadata$meter_index <= runtime_meter_idx;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_storm_control_meter_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetStormControlMeterRspT {pkt: pkt, meter_metadata$meter_index: meter_metadata$meter_index};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_STP_STATE ======

interface SetStpState;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetStpState  (SetStpState);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$stp_state <- mkReg(0);
  rule set_stp_state_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetStpStateReqT {pkt: .pkt, runtime_stp_state: .runtime_stp_state}: begin
        l2_metadata$stp_state <= runtime_stp_state;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_stp_state_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetStpStateRspT {pkt: pkt, l2_metadata$stp_state: l2_metadata$stp_state};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_TUNNEL_REWRITE_DETAILS ======

interface SetTunnelRewriteDetails;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetTunnelRewriteDetails  (SetTunnelRewriteDetails);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) egress_metadata$outer_bd <- mkReg(0);
  Reg#(Bit#(9)) tunnel_metadata$tunnel_smac_index <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_dmac_index <- mkReg(0);
  Reg#(Bit#(9)) tunnel_metadata$tunnel_src_index <- mkReg(0);
  Reg#(Bit#(14)) tunnel_metadata$tunnel_dst_index <- mkReg(0);
  rule set_tunnel_rewrite_details_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetTunnelRewriteDetailsReqT {pkt: .pkt, runtime_outer_bd: .runtime_outer_bd, runtime_sip_index: .runtime_sip_index, runtime_dip_index: .runtime_dip_index, runtime_dmac_idx: .runtime_dmac_idx, runtime_smac_idx: .runtime_smac_idx}: begin
        egress_metadata$outer_bd <= runtime_outer_bd;
        tunnel_metadata$tunnel_smac_index <= runtime_smac_idx;
        tunnel_metadata$tunnel_dmac_index <= runtime_dmac_idx;
        tunnel_metadata$tunnel_src_index <= runtime_sip_index;
        tunnel_metadata$tunnel_dst_index <= runtime_dip_index;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_tunnel_rewrite_details_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetTunnelRewriteDetailsRspT {pkt: pkt, egress_metadata$outer_bd: egress_metadata$outer_bd, tunnel_metadata$tunnel_src_index: tunnel_metadata$tunnel_src_index, tunnel_metadata$tunnel_dst_index: tunnel_metadata$tunnel_dst_index, tunnel_metadata$tunnel_dmac_index: tunnel_metadata$tunnel_dmac_index, tunnel_metadata$tunnel_smac_index: tunnel_metadata$tunnel_smac_index};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_TUNNEL_TERMINATION_FLAG ======

interface SetTunnelTerminationFlag;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetTunnelTerminationFlag  (SetTunnelTerminationFlag);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  rule set_tunnel_termination_flag_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetTunnelTerminationFlagReqT {pkt: .pkt}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_tunnel_termination_flag_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetTunnelTerminationFlagRspT {pkt: pkt, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_TUNNEL_VNI_AND_TERMINATION_FLAG ======

interface SetTunnelVniAndTerminationFlag;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetTunnelVniAndTerminationFlag  (SetTunnelVniAndTerminationFlag);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(24)) tunnel_metadata$tunnel_vni <- mkReg(0);
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  rule set_tunnel_vni_and_termination_flag_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetTunnelVniAndTerminationFlagReqT {pkt: .pkt, runtime_tunnel_vni: .runtime_tunnel_vni}: begin
        tunnel_metadata$tunnel_vni <= runtime_tunnel_vni;
        tunnel_metadata$tunnel_terminate <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_tunnel_vni_and_termination_flag_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetTunnelVniAndTerminationFlagRspT {pkt: pkt, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, tunnel_metadata$tunnel_vni: tunnel_metadata$tunnel_vni};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_UNICAST ======

interface SetUnicast;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetUnicast  (SetUnicast);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  rule set_unicast_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetUnicastReqT {pkt: .pkt}: begin
        l2_metadata$lkp_pkt_type <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_unicast_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetUnicastRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_UNICAST_AND_IPV6_SRC_IS_LINK_LOCAL ======

interface SetUnicastAndIpv6SrcIsLinkLocal;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetUnicastAndIpv6SrcIsLinkLocal  (SetUnicastAndIpv6SrcIsLinkLocal);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(1)) ipv6_metadata$ipv6_src_is_link_local <- mkReg(0);
  rule set_unicast_and_ipv6_src_is_link_local_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetUnicastAndIpv6SrcIsLinkLocalReqT {pkt: .pkt}: begin
        l2_metadata$lkp_pkt_type <= 'h1;
        ipv6_metadata$ipv6_src_is_link_local <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_unicast_and_ipv6_src_is_link_local_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetUnicastAndIpv6SrcIsLinkLocalRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, ipv6_metadata$ipv6_src_is_link_local: ipv6_metadata$ipv6_src_is_link_local};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_MPLS_LABEL1 ======

interface SetValidMplsLabel1;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidMplsLabel1  (SetValidMplsLabel1);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(20)) tunnel_metadata$mpls_label <- mkReg(0);
  Reg#(Bit#(3)) tunnel_metadata$mpls_exp <- mkReg(0);
  rule set_valid_mpls_label1_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidMplsLabel1ReqT {pkt: .pkt, mpls0$exp: .mpls0$exp, mpls0$label: .mpls0$label}: begin
        tunnel_metadata$mpls_label <= mpls0$label;
        tunnel_metadata$mpls_exp <= mpls0$exp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_mpls_label1_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidMplsLabel1RspT {pkt: pkt, tunnel_metadata$mpls_label: tunnel_metadata$mpls_label, tunnel_metadata$mpls_exp: tunnel_metadata$mpls_exp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_MPLS_LABEL2 ======

interface SetValidMplsLabel2;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidMplsLabel2  (SetValidMplsLabel2);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(20)) tunnel_metadata$mpls_label <- mkReg(0);
  Reg#(Bit#(3)) tunnel_metadata$mpls_exp <- mkReg(0);
  rule set_valid_mpls_label2_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidMplsLabel2ReqT {pkt: .pkt, mpls1$label: .mpls1$label, mpls1$exp: .mpls1$exp}: begin
        tunnel_metadata$mpls_label <= mpls1$label;
        tunnel_metadata$mpls_exp <= mpls1$exp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_mpls_label2_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidMplsLabel2RspT {pkt: pkt, tunnel_metadata$mpls_label: tunnel_metadata$mpls_label, tunnel_metadata$mpls_exp: tunnel_metadata$mpls_exp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_MPLS_LABEL3 ======

interface SetValidMplsLabel3;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidMplsLabel3  (SetValidMplsLabel3);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(20)) tunnel_metadata$mpls_label <- mkReg(0);
  Reg#(Bit#(3)) tunnel_metadata$mpls_exp <- mkReg(0);
  rule set_valid_mpls_label3_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidMplsLabel3ReqT {pkt: .pkt, mpls2$label: .mpls2$label, mpls2$exp: .mpls2$exp}: begin
        tunnel_metadata$mpls_label <= mpls2$label;
        tunnel_metadata$mpls_exp <= mpls2$exp;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_mpls_label3_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidMplsLabel3RspT {pkt: pkt, tunnel_metadata$mpls_label: tunnel_metadata$mpls_label, tunnel_metadata$mpls_exp: tunnel_metadata$mpls_exp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_BROADCAST_PACKET_DOUBLE_TAGGED ======

interface SetValidOuterBroadcastPacketDoubleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterBroadcastPacketDoubleTagged  (SetValidOuterBroadcastPacketDoubleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_broadcast_packet_double_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterBroadcastPacketDoubleTaggedReqT {pkt: .pkt, vlan_tag_1$etherType: .vlan_tag_1$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h4;
        l2_metadata$lkp_mac_type <= vlan_tag_1$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_broadcast_packet_double_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterBroadcastPacketDoubleTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_BROADCAST_PACKET_QINQ_TAGGED ======

interface SetValidOuterBroadcastPacketQinqTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterBroadcastPacketQinqTagged  (SetValidOuterBroadcastPacketQinqTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_broadcast_packet_qinq_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterBroadcastPacketQinqTaggedReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h4;
        l2_metadata$lkp_mac_type <= ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_broadcast_packet_qinq_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterBroadcastPacketQinqTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_BROADCAST_PACKET_SINGLE_TAGGED ======

interface SetValidOuterBroadcastPacketSingleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterBroadcastPacketSingleTagged  (SetValidOuterBroadcastPacketSingleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_broadcast_packet_single_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterBroadcastPacketSingleTaggedReqT {pkt: .pkt, vlan_tag_0$etherType: .vlan_tag_0$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h4;
        l2_metadata$lkp_mac_type <= vlan_tag_0$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_broadcast_packet_single_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterBroadcastPacketSingleTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_BROADCAST_PACKET_UNTAGGED ======

interface SetValidOuterBroadcastPacketUntagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterBroadcastPacketUntagged  (SetValidOuterBroadcastPacketUntagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_broadcast_packet_untagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterBroadcastPacketUntaggedReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h4;
        l2_metadata$lkp_mac_type <= ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_broadcast_packet_untagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterBroadcastPacketUntaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_IPV4_PACKET ======

interface SetValidOuterIpv4Packet;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterIpv4Packet  (SetValidOuterIpv4Packet);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_tc <- mkReg(0);
  Reg#(Bit#(4)) l3_metadata$lkp_ip_version <- mkReg(0);
  rule set_valid_outer_ipv4_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterIpv4PacketReqT {pkt: .pkt, ipv4$diffserv: .ipv4$diffserv, ipv4$version: .ipv4$version}: begin
        l3_metadata$lkp_ip_type <= 'h1;
        l3_metadata$lkp_ip_tc <= ipv4$diffserv;
        l3_metadata$lkp_ip_version <= ipv4$version;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_ipv4_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterIpv4PacketRspT {pkt: pkt, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_IPV6_PACKET ======

interface SetValidOuterIpv6Packet;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterIpv6Packet  (SetValidOuterIpv6Packet);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_tc <- mkReg(0);
  Reg#(Bit#(4)) l3_metadata$lkp_ip_version <- mkReg(0);
  rule set_valid_outer_ipv6_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterIpv6PacketReqT {pkt: .pkt, ipv6$version: .ipv6$version, ipv6$trafficClass: .ipv6$trafficClass}: begin
        l3_metadata$lkp_ip_type <= 'h2;
        l3_metadata$lkp_ip_tc <= ipv6$trafficClass;
        l3_metadata$lkp_ip_version <= ipv6$version;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_ipv6_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterIpv6PacketRspT {pkt: pkt, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_MULTICAST_PACKET_DOUBLE_TAGGED ======

interface SetValidOuterMulticastPacketDoubleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterMulticastPacketDoubleTagged  (SetValidOuterMulticastPacketDoubleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_multicast_packet_double_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterMulticastPacketDoubleTaggedReqT {pkt: .pkt, vlan_tag_1$etherType: .vlan_tag_1$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h2;
        l2_metadata$lkp_mac_type <= vlan_tag_1$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_multicast_packet_double_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterMulticastPacketDoubleTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_MULTICAST_PACKET_QINQ_TAGGED ======

interface SetValidOuterMulticastPacketQinqTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterMulticastPacketQinqTagged  (SetValidOuterMulticastPacketQinqTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_multicast_packet_qinq_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterMulticastPacketQinqTaggedReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h2;
        l2_metadata$lkp_mac_type <= ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_multicast_packet_qinq_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterMulticastPacketQinqTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_MULTICAST_PACKET_SINGLE_TAGGED ======

interface SetValidOuterMulticastPacketSingleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterMulticastPacketSingleTagged  (SetValidOuterMulticastPacketSingleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_multicast_packet_single_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterMulticastPacketSingleTaggedReqT {pkt: .pkt, vlan_tag_0$etherType: .vlan_tag_0$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h2;
        l2_metadata$lkp_mac_type <= vlan_tag_0$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_multicast_packet_single_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterMulticastPacketSingleTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_MULTICAST_PACKET_UNTAGGED ======

interface SetValidOuterMulticastPacketUntagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterMulticastPacketUntagged  (SetValidOuterMulticastPacketUntagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_multicast_packet_untagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterMulticastPacketUntaggedReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h2;
        l2_metadata$lkp_mac_type <= ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_multicast_packet_untagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterMulticastPacketUntaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_UNICAST_PACKET_DOUBLE_TAGGED ======

interface SetValidOuterUnicastPacketDoubleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterUnicastPacketDoubleTagged  (SetValidOuterUnicastPacketDoubleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_unicast_packet_double_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterUnicastPacketDoubleTaggedReqT {pkt: .pkt, vlan_tag_1$etherType: .vlan_tag_1$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h1;
        l2_metadata$lkp_mac_type <= vlan_tag_1$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_unicast_packet_double_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterUnicastPacketDoubleTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_UNICAST_PACKET_QINQ_TAGGED ======

interface SetValidOuterUnicastPacketQinqTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterUnicastPacketQinqTagged  (SetValidOuterUnicastPacketQinqTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_unicast_packet_qinq_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterUnicastPacketQinqTaggedReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h1;
        l2_metadata$lkp_mac_type <= ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_unicast_packet_qinq_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterUnicastPacketQinqTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_UNICAST_PACKET_SINGLE_TAGGED ======

interface SetValidOuterUnicastPacketSingleTagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterUnicastPacketSingleTagged  (SetValidOuterUnicastPacketSingleTagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_unicast_packet_single_tagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterUnicastPacketSingleTaggedReqT {pkt: .pkt, vlan_tag_0$etherType: .vlan_tag_0$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h1;
        l2_metadata$lkp_mac_type <= vlan_tag_0$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_unicast_packet_single_tagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterUnicastPacketSingleTaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SET_VALID_OUTER_UNICAST_PACKET_UNTAGGED ======

interface SetValidOuterUnicastPacketUntagged;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSetValidOuterUnicastPacketUntagged  (SetValidOuterUnicastPacketUntagged);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(3)) l2_metadata$lkp_pkt_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule set_valid_outer_unicast_packet_untagged_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SetValidOuterUnicastPacketUntaggedReqT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        l2_metadata$lkp_pkt_type <= 'h1;
        l2_metadata$lkp_mac_type <= ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule set_valid_outer_unicast_packet_untagged_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SetValidOuterUnicastPacketUntaggedRspT {pkt: pkt, l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SFLOW_ING_PKT_TO_CPU ======

interface SflowIngPktToCpu;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSflowIngPktToCpu  (SflowIngPktToCpu);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) fabric_metadata$reason_code <- mkReg(0);
  Reg#(Bit#(16)) i2e_metadata$mirror_session_id <- mkReg(0);
  rule sflow_ing_pkt_to_cpu_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SflowIngPktToCpuReqT {pkt: .pkt, runtime_sflow_i2e_mirror_id: .runtime_sflow_i2e_mirror_id, runtime_reason_code: .runtime_reason_code}: begin
        fabric_metadata$reason_code <= runtime_reason_code;
        i2e_metadata$mirror_session_id <= runtime_sflow_i2e_mirror_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule sflow_ing_pkt_to_cpu_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SflowIngPktToCpuRspT {pkt: pkt, fabric_metadata$reason_code: fabric_metadata$reason_code, i2e_metadata$mirror_session_id: i2e_metadata$mirror_session_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SFLOW_ING_SESSION_ENABLE ======

interface SflowIngSessionEnable;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSflowIngSessionEnable  (SflowIngSessionEnable);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) sflow_metadata$sflow_session_id <- mkReg(0);
  rule sflow_ing_session_enable_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SflowIngSessionEnableReqT {pkt: .pkt, runtime_rate_thr: .runtime_rate_thr, runtime_session_id: .runtime_session_id}: begin
        sflow_metadata$sflow_session_id <= runtime_session_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule sflow_ing_session_enable_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SflowIngSessionEnableRspT {pkt: pkt, sflow_metadata$sflow_session_id: sflow_metadata$sflow_session_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SFLOW_PKT_TO_CPU ======

interface SflowPktToCpu;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSflowPktToCpu  (SflowPktToCpu);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) fabric_header_sflow$sflow_session_id <- mkReg(0);
  rule sflow_pkt_to_cpu_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SflowPktToCpuReqT {pkt: .pkt, sflow_metadata$sflow_session_id: .sflow_metadata$sflow_session_id}: begin
        fabric_header_sflow$sflow_session_id <= sflow_metadata$sflow_session_id;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule sflow_pkt_to_cpu_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SflowPktToCpuRspT {pkt: pkt, fabric_header_sflow$sflow_session_id: fabric_header_sflow$sflow_session_id};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SMAC_HIT ======

interface SmacHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSmacHit  (SmacHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule smac_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SmacHitReqT {pkt: .pkt, runtime_ifindex: .runtime_ifindex}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule smac_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SmacHitRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SMAC_MISS ======

interface SmacMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSmacMiss  (SmacMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l2_metadata$l2_src_miss <- mkReg(0);
  rule smac_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SmacMissReqT {pkt: .pkt}: begin
        l2_metadata$l2_src_miss <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule smac_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SmacMissRspT {pkt: pkt, l2_metadata$l2_src_miss: l2_metadata$l2_src_miss};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SRC_VTEP_HIT ======

interface SrcVtepHit;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSrcVtepHit  (SrcVtepHit);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ingress_metadata$ifindex <- mkReg(0);
  rule src_vtep_hit_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SrcVtepHitReqT {pkt: .pkt, runtime_ifindex: .runtime_ifindex}: begin
        ingress_metadata$ifindex <= runtime_ifindex;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule src_vtep_hit_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SrcVtepHitRspT {pkt: pkt, ingress_metadata$ifindex: ingress_metadata$ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SWITCH_FABRIC_MULTICAST_PACKET ======

interface SwitchFabricMulticastPacket;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSwitchFabricMulticastPacket  (SwitchFabricMulticastPacket);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) fabric_metadata$fabric_header_present <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  rule switch_fabric_multicast_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SwitchFabricMulticastPacketReqT {pkt: .pkt, fabric_header$dstPortOrGroup: .fabric_header$dstPortOrGroup}: begin
        fabric_metadata$fabric_header_present <= 'h1;
        intrinsic_metadata$mcast_grp <= fabric_header$dstPortOrGroup;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule switch_fabric_multicast_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SwitchFabricMulticastPacketRspT {pkt: pkt, fabric_metadata$fabric_header_present: fabric_metadata$fabric_header_present, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== SWITCH_FABRIC_UNICAST_PACKET ======

interface SwitchFabricUnicastPacket;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkSwitchFabricUnicastPacket  (SwitchFabricUnicastPacket);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) fabric_metadata$fabric_header_present <- mkReg(0);
  Reg#(Bit#(8)) fabric_metadata$dst_device <- mkReg(0);
  Reg#(Bit#(16)) fabric_metadata$dst_port <- mkReg(0);
  rule switch_fabric_unicast_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged SwitchFabricUnicastPacketReqT {pkt: .pkt, fabric_header$dstDevice: .fabric_header$dstDevice, fabric_header$dstPortOrGroup: .fabric_header$dstPortOrGroup}: begin
        fabric_metadata$fabric_header_present <= 'h1;
        fabric_metadata$dst_device <= fabric_header$dstDevice;
        fabric_metadata$dst_port <= fabric_header$dstPortOrGroup;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule switch_fabric_unicast_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged SwitchFabricUnicastPacketRspT {pkt: pkt, fabric_metadata$fabric_header_present: fabric_metadata$fabric_header_present, fabric_metadata$dst_port: fabric_metadata$dst_port, fabric_metadata$dst_device: fabric_metadata$dst_device};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_CPU_PACKET ======

interface TerminateCpuPacket;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateCpuPacket  (TerminateCpuPacket);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(9)) standard_metadata$egress_spec <- mkReg(0);
  Reg#(Bit#(1)) egress_metadata$bypass <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule terminate_cpu_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateCpuPacketReqT {pkt: .pkt, fabric_payload_header$etherType: .fabric_payload_header$etherType, fabric_header_cpu$txBypass: .fabric_header_cpu$txBypass, fabric_header$dstPortOrGroup: .fabric_header$dstPortOrGroup}: begin
        standard_metadata$egress_spec <= fabric_header$dstPortOrGroup;
        egress_metadata$bypass <= fabric_header_cpu$txBypass;
        ethernet$etherType <= fabric_payload_header$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_cpu_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateCpuPacketRspT {pkt: pkt, egress_metadata$bypass: egress_metadata$bypass, standard_metadata$egress_spec: standard_metadata$egress_spec, ethernet$etherType: ethernet$etherType};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_EOMPLS ======

interface TerminateEompls;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateEompls  (TerminateEompls);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$ingress_tunnel_type <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule terminate_eompls_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateEomplsReqT {pkt: .pkt, inner_ethernet$etherType: .inner_ethernet$etherType, runtime_tunnel_type: .runtime_tunnel_type, runtime_bd: .runtime_bd}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        tunnel_metadata$ingress_tunnel_type <= runtime_tunnel_type;
        ingress_metadata$bd <= runtime_bd;
        l2_metadata$lkp_mac_type <= inner_ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_eompls_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateEomplsRspT {pkt: pkt, tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type, ingress_metadata$bd: ingress_metadata$bd};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_FABRIC_MULTICAST_PACKET ======

interface TerminateFabricMulticastPacket;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateFabricMulticastPacket  (TerminateFabricMulticastPacket);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$ingress_tunnel_type <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$routed <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$outer_routed <- mkReg(0);
  Reg#(Bit#(16)) intrinsic_metadata$mcast_grp <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule terminate_fabric_multicast_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateFabricMulticastPacketReqT {pkt: .pkt, fabric_payload_header$etherType: .fabric_payload_header$etherType, fabric_header_multicast$tunnelTerminate: .fabric_header_multicast$tunnelTerminate, fabric_header_multicast$outerRouted: .fabric_header_multicast$outerRouted, fabric_header_multicast$ingressTunnelType: .fabric_header_multicast$ingressTunnelType, fabric_header_multicast$mcastGrp: .fabric_header_multicast$mcastGrp, fabric_header_multicast$routed: .fabric_header_multicast$routed}: begin
        tunnel_metadata$tunnel_terminate <= fabric_header_multicast$tunnelTerminate;
        tunnel_metadata$ingress_tunnel_type <= fabric_header_multicast$ingressTunnelType;
        l3_metadata$nexthop_index <= 'h0;
        l3_metadata$routed <= fabric_header_multicast$routed;
        l3_metadata$outer_routed <= fabric_header_multicast$outerRouted;
        intrinsic_metadata$mcast_grp <= fabric_header_multicast$mcastGrp;
        ethernet$etherType <= fabric_payload_header$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_fabric_multicast_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateFabricMulticastPacketRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp, l3_metadata$routed: l3_metadata$routed, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, ethernet$etherType: ethernet$etherType, l3_metadata$outer_routed: l3_metadata$outer_routed};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_FABRIC_UNICAST_PACKET ======

interface TerminateFabricUnicastPacket;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateFabricUnicastPacket  (TerminateFabricUnicastPacket);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(9)) standard_metadata$egress_spec <- mkReg(0);
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$ingress_tunnel_type <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$nexthop_index <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$routed <- mkReg(0);
  Reg#(Bit#(1)) l3_metadata$outer_routed <- mkReg(0);
  Reg#(Bit#(16)) ethernet$etherType <- mkReg(0);
  rule terminate_fabric_unicast_packet_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateFabricUnicastPacketReqT {pkt: .pkt, fabric_header_unicast$nexthopIndex: .fabric_header_unicast$nexthopIndex, fabric_header_unicast$routed: .fabric_header_unicast$routed, fabric_header_unicast$tunnelTerminate: .fabric_header_unicast$tunnelTerminate, fabric_payload_header$etherType: .fabric_payload_header$etherType, fabric_header_unicast$outerRouted: .fabric_header_unicast$outerRouted, fabric_header_unicast$ingressTunnelType: .fabric_header_unicast$ingressTunnelType, fabric_header$dstPortOrGroup: .fabric_header$dstPortOrGroup}: begin
        standard_metadata$egress_spec <= fabric_header$dstPortOrGroup;
        tunnel_metadata$tunnel_terminate <= fabric_header_unicast$tunnelTerminate;
        tunnel_metadata$ingress_tunnel_type <= fabric_header_unicast$ingressTunnelType;
        l3_metadata$nexthop_index <= fabric_header_unicast$nexthopIndex;
        l3_metadata$routed <= fabric_header_unicast$routed;
        l3_metadata$outer_routed <= fabric_header_unicast$outerRouted;
        ethernet$etherType <= fabric_payload_header$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_fabric_unicast_packet_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateFabricUnicastPacketRspT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type, standard_metadata$egress_spec: standard_metadata$egress_spec, l3_metadata$routed: l3_metadata$routed, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, ethernet$etherType: ethernet$etherType, l3_metadata$outer_routed: l3_metadata$outer_routed};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_IPV4_OVER_MPLS ======

interface TerminateIpv4OverMpls;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateIpv4OverMpls  (TerminateIpv4OverMpls);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$ingress_tunnel_type <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$vrf <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  Reg#(Bit#(4)) l3_metadata$lkp_ip_version <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_tc <- mkReg(0);
  rule terminate_ipv4_over_mpls_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateIpv4OverMplsReqT {pkt: .pkt, inner_ipv4$diffserv: .inner_ipv4$diffserv, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, inner_ethernet$etherType: .inner_ethernet$etherType, inner_ipv4$version: .inner_ipv4$version, runtime_tunnel_type: .runtime_tunnel_type, runtime_vrf: .runtime_vrf}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        tunnel_metadata$ingress_tunnel_type <= runtime_tunnel_type;
        l3_metadata$vrf <= runtime_vrf;
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        l3_metadata$lkp_ip_type <= 'h1;
        l2_metadata$lkp_mac_type <= inner_ethernet$etherType;
        l3_metadata$lkp_ip_version <= inner_ipv4$version;
        l3_metadata$lkp_ip_tc <= inner_ipv4$diffserv;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_ipv4_over_mpls_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateIpv4OverMplsRspT {pkt: pkt, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, l3_metadata$vrf: l3_metadata$vrf, l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_IPV6_OVER_MPLS ======

interface TerminateIpv6OverMpls;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateIpv6OverMpls  (TerminateIpv6OverMpls);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$ingress_tunnel_type <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$vrf <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  Reg#(Bit#(4)) l3_metadata$lkp_ip_version <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_tc <- mkReg(0);
  rule terminate_ipv6_over_mpls_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateIpv6OverMplsReqT {pkt: .pkt, inner_ipv6$version: .inner_ipv6$version, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, inner_ethernet$etherType: .inner_ethernet$etherType, inner_ipv6$trafficClass: .inner_ipv6$trafficClass, runtime_tunnel_type: .runtime_tunnel_type, runtime_vrf: .runtime_vrf}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        tunnel_metadata$ingress_tunnel_type <= runtime_tunnel_type;
        l3_metadata$vrf <= runtime_vrf;
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        l3_metadata$lkp_ip_type <= 'h2;
        l2_metadata$lkp_mac_type <= inner_ethernet$etherType;
        l3_metadata$lkp_ip_version <= inner_ipv6$version;
        l3_metadata$lkp_ip_tc <= inner_ipv6$trafficClass;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_ipv6_over_mpls_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateIpv6OverMplsRspT {pkt: pkt, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, l3_metadata$vrf: l3_metadata$vrf, l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_PW ======

interface TerminatePw;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminatePw  (TerminatePw);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) ingress_metadata$egress_ifindex <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  rule terminate_pw_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminatePwReqT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, runtime_ifindex: .runtime_ifindex}: begin
        ingress_metadata$egress_ifindex <= runtime_ifindex;
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_pw_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminatePwRspT {pkt: pkt, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da, ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_TUNNEL_INNER_ETHERNET_IPV4 ======

interface TerminateTunnelInnerEthernetIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateTunnelInnerEthernetIpv4  (TerminateTunnelInnerEthernetIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$vrf <- mkReg(0);
  Reg#(Bit#(8)) qos_metadata$outer_dscp <- mkReg(0);
  Reg#(Bit#(1)) ipv4_metadata$ipv4_unicast_enabled <- mkReg(0);
  Reg#(Bit#(2)) ipv4_metadata$ipv4_urpf_mode <- mkReg(0);
  Reg#(Bit#(10)) l3_metadata$rmac_group <- mkReg(0);
  Reg#(Bit#(16)) acl_metadata$bd_label <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$bd_stats_idx <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  Reg#(Bit#(4)) l3_metadata$lkp_ip_version <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_tc <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$igmp_snooping_enabled <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$ipv4_multicast_enabled <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$bd_mrpf_group <- mkReg(0);
  rule terminate_tunnel_inner_ethernet_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateTunnelInnerEthernetIpv4ReqT {pkt: .pkt, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, inner_ipv4$version: .inner_ipv4$version, inner_ethernet$etherType: .inner_ethernet$etherType, inner_ipv4$diffserv: .inner_ipv4$diffserv, runtime_ipv4_multicast_enabled: .runtime_ipv4_multicast_enabled, runtime_igmp_snooping_enabled: .runtime_igmp_snooping_enabled, runtime_mrpf_group: .runtime_mrpf_group, runtime_stats_idx: .runtime_stats_idx, runtime_ipv4_urpf_mode: .runtime_ipv4_urpf_mode, runtime_bd: .runtime_bd, runtime_vrf: .runtime_vrf, runtime_bd_label: .runtime_bd_label, runtime_rmac_group: .runtime_rmac_group, runtime_ipv4_unicast_enabled: .runtime_ipv4_unicast_enabled}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        ingress_metadata$bd <= runtime_bd;
        l3_metadata$vrf <= runtime_vrf;
        qos_metadata$outer_dscp <= l3_metadata$lkp_ip_tc;
        ipv4_metadata$ipv4_unicast_enabled <= runtime_ipv4_unicast_enabled;
        ipv4_metadata$ipv4_urpf_mode <= runtime_ipv4_urpf_mode;
        l3_metadata$rmac_group <= runtime_rmac_group;
        acl_metadata$bd_label <= runtime_bd_label;
        l2_metadata$bd_stats_idx <= runtime_stats_idx;
        l3_metadata$lkp_ip_type <= 'h1;
        l2_metadata$lkp_mac_type <= inner_ethernet$etherType;
        l3_metadata$lkp_ip_version <= inner_ipv4$version;
        l3_metadata$lkp_ip_tc <= inner_ipv4$diffserv;
        multicast_metadata$igmp_snooping_enabled <= runtime_igmp_snooping_enabled;
        multicast_metadata$ipv4_multicast_enabled <= runtime_ipv4_multicast_enabled;
        multicast_metadata$bd_mrpf_group <= runtime_mrpf_group;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_tunnel_inner_ethernet_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateTunnelInnerEthernetIpv4RspT {pkt: pkt, l3_metadata$rmac_group: l3_metadata$rmac_group, multicast_metadata$igmp_snooping_enabled: multicast_metadata$igmp_snooping_enabled, multicast_metadata$bd_mrpf_group: multicast_metadata$bd_mrpf_group, multicast_metadata$ipv4_multicast_enabled: multicast_metadata$ipv4_multicast_enabled, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type, acl_metadata$bd_label: acl_metadata$bd_label, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, l3_metadata$vrf: l3_metadata$vrf, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version, qos_metadata$outer_dscp: qos_metadata$outer_dscp, ingress_metadata$bd: ingress_metadata$bd, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, ipv4_metadata$ipv4_urpf_mode: ipv4_metadata$ipv4_urpf_mode, l2_metadata$bd_stats_idx: l2_metadata$bd_stats_idx, ipv4_metadata$ipv4_unicast_enabled: ipv4_metadata$ipv4_unicast_enabled};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_TUNNEL_INNER_ETHERNET_IPV6 ======

interface TerminateTunnelInnerEthernetIpv6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateTunnelInnerEthernetIpv6  (TerminateTunnelInnerEthernetIpv6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$vrf <- mkReg(0);
  Reg#(Bit#(8)) qos_metadata$outer_dscp <- mkReg(0);
  Reg#(Bit#(1)) ipv6_metadata$ipv6_unicast_enabled <- mkReg(0);
  Reg#(Bit#(2)) ipv6_metadata$ipv6_urpf_mode <- mkReg(0);
  Reg#(Bit#(10)) l3_metadata$rmac_group <- mkReg(0);
  Reg#(Bit#(16)) acl_metadata$bd_label <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$bd_stats_idx <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  Reg#(Bit#(4)) l3_metadata$lkp_ip_version <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_tc <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$bd_mrpf_group <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$ipv6_multicast_enabled <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$mld_snooping_enabled <- mkReg(0);
  rule terminate_tunnel_inner_ethernet_ipv6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateTunnelInnerEthernetIpv6ReqT {pkt: .pkt, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, inner_ipv6$trafficClass: .inner_ipv6$trafficClass, inner_ethernet$etherType: .inner_ethernet$etherType, inner_ipv6$version: .inner_ipv6$version, runtime_mrpf_group: .runtime_mrpf_group, runtime_mld_snooping_enabled: .runtime_mld_snooping_enabled, runtime_ipv6_multicast_enabled: .runtime_ipv6_multicast_enabled, runtime_stats_idx: .runtime_stats_idx, runtime_ipv6_urpf_mode: .runtime_ipv6_urpf_mode, runtime_bd: .runtime_bd, runtime_vrf: .runtime_vrf, runtime_ipv6_unicast_enabled: .runtime_ipv6_unicast_enabled, runtime_bd_label: .runtime_bd_label, runtime_rmac_group: .runtime_rmac_group}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        ingress_metadata$bd <= runtime_bd;
        l3_metadata$vrf <= runtime_vrf;
        qos_metadata$outer_dscp <= l3_metadata$lkp_ip_tc;
        ipv6_metadata$ipv6_unicast_enabled <= runtime_ipv6_unicast_enabled;
        ipv6_metadata$ipv6_urpf_mode <= runtime_ipv6_urpf_mode;
        l3_metadata$rmac_group <= runtime_rmac_group;
        acl_metadata$bd_label <= runtime_bd_label;
        l2_metadata$bd_stats_idx <= runtime_stats_idx;
        l3_metadata$lkp_ip_type <= 'h2;
        l2_metadata$lkp_mac_type <= inner_ethernet$etherType;
        l3_metadata$lkp_ip_version <= inner_ipv6$version;
        l3_metadata$lkp_ip_tc <= inner_ipv6$trafficClass;
        multicast_metadata$bd_mrpf_group <= runtime_mrpf_group;
        multicast_metadata$ipv6_multicast_enabled <= runtime_ipv6_multicast_enabled;
        multicast_metadata$mld_snooping_enabled <= runtime_mld_snooping_enabled;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_tunnel_inner_ethernet_ipv6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateTunnelInnerEthernetIpv6RspT {pkt: pkt, l3_metadata$rmac_group: l3_metadata$rmac_group, multicast_metadata$bd_mrpf_group: multicast_metadata$bd_mrpf_group, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type, acl_metadata$bd_label: acl_metadata$bd_label, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, l3_metadata$vrf: l3_metadata$vrf, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, ipv6_metadata$ipv6_unicast_enabled: ipv6_metadata$ipv6_unicast_enabled, ipv6_metadata$ipv6_urpf_mode: ipv6_metadata$ipv6_urpf_mode, qos_metadata$outer_dscp: qos_metadata$outer_dscp, ingress_metadata$bd: ingress_metadata$bd, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, multicast_metadata$ipv6_multicast_enabled: multicast_metadata$ipv6_multicast_enabled, l2_metadata$bd_stats_idx: l2_metadata$bd_stats_idx, l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version, multicast_metadata$mld_snooping_enabled: multicast_metadata$mld_snooping_enabled};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_TUNNEL_INNER_IPV4 ======

interface TerminateTunnelInnerIpv4;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateTunnelInnerIpv4  (TerminateTunnelInnerIpv4);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$vrf <- mkReg(0);
  Reg#(Bit#(8)) qos_metadata$outer_dscp <- mkReg(0);
  Reg#(Bit#(1)) ipv4_metadata$ipv4_unicast_enabled <- mkReg(0);
  Reg#(Bit#(2)) ipv4_metadata$ipv4_urpf_mode <- mkReg(0);
  Reg#(Bit#(10)) l3_metadata$rmac_group <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(4)) l3_metadata$lkp_ip_version <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_tc <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$bd_mrpf_group <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$ipv4_multicast_enabled <- mkReg(0);
  rule terminate_tunnel_inner_ipv4_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateTunnelInnerIpv4ReqT {pkt: .pkt, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, inner_ipv4$diffserv: .inner_ipv4$diffserv, inner_ipv4$version: .inner_ipv4$version, runtime_ipv4_multicast_enabled: .runtime_ipv4_multicast_enabled, runtime_mrpf_group: .runtime_mrpf_group, runtime_ipv4_urpf_mode: .runtime_ipv4_urpf_mode, runtime_vrf: .runtime_vrf, runtime_rmac_group: .runtime_rmac_group, runtime_ipv4_unicast_enabled: .runtime_ipv4_unicast_enabled}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        l3_metadata$vrf <= runtime_vrf;
        qos_metadata$outer_dscp <= l3_metadata$lkp_ip_tc;
        ipv4_metadata$ipv4_unicast_enabled <= runtime_ipv4_unicast_enabled;
        ipv4_metadata$ipv4_urpf_mode <= runtime_ipv4_urpf_mode;
        l3_metadata$rmac_group <= runtime_rmac_group;
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        l3_metadata$lkp_ip_type <= 'h1;
        l3_metadata$lkp_ip_version <= inner_ipv4$version;
        l3_metadata$lkp_ip_tc <= inner_ipv4$diffserv;
        multicast_metadata$bd_mrpf_group <= runtime_mrpf_group;
        multicast_metadata$ipv4_multicast_enabled <= runtime_ipv4_multicast_enabled;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_tunnel_inner_ipv4_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateTunnelInnerIpv4RspT {pkt: pkt, l3_metadata$rmac_group: l3_metadata$rmac_group, ipv4_metadata$ipv4_urpf_mode: ipv4_metadata$ipv4_urpf_mode, multicast_metadata$bd_mrpf_group: multicast_metadata$bd_mrpf_group, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, l3_metadata$vrf: l3_metadata$vrf, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, multicast_metadata$ipv4_multicast_enabled: multicast_metadata$ipv4_multicast_enabled, qos_metadata$outer_dscp: qos_metadata$outer_dscp, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, ipv4_metadata$ipv4_unicast_enabled: ipv4_metadata$ipv4_unicast_enabled, l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_TUNNEL_INNER_IPV6 ======

interface TerminateTunnelInnerIpv6;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateTunnelInnerIpv6  (TerminateTunnelInnerIpv6);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(16)) l3_metadata$vrf <- mkReg(0);
  Reg#(Bit#(8)) qos_metadata$outer_dscp <- mkReg(0);
  Reg#(Bit#(1)) ipv6_metadata$ipv6_unicast_enabled <- mkReg(0);
  Reg#(Bit#(2)) ipv6_metadata$ipv6_urpf_mode <- mkReg(0);
  Reg#(Bit#(10)) l3_metadata$rmac_group <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_sa <- mkReg(0);
  Reg#(Bit#(48)) l2_metadata$lkp_mac_da <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(128)) ipv6_metadata$lkp_ipv6_sa <- mkReg(0);
  Reg#(Bit#(128)) ipv6_metadata$lkp_ipv6_da <- mkReg(0);
  Reg#(Bit#(4)) l3_metadata$lkp_ip_version <- mkReg(0);
  Reg#(Bit#(8)) l3_metadata$lkp_ip_tc <- mkReg(0);
  Reg#(Bit#(16)) multicast_metadata$bd_mrpf_group <- mkReg(0);
  Reg#(Bit#(1)) multicast_metadata$ipv6_multicast_enabled <- mkReg(0);
  rule terminate_tunnel_inner_ipv6_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateTunnelInnerIpv6ReqT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr, ethernet$dstAddr: .ethernet$dstAddr, inner_ipv6$dstAddr: .inner_ipv6$dstAddr, inner_ipv6$srcAddr: .inner_ipv6$srcAddr, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, inner_ipv6$trafficClass: .inner_ipv6$trafficClass, inner_ipv6$version: .inner_ipv6$version, runtime_mrpf_group: .runtime_mrpf_group, runtime_ipv6_multicast_enabled: .runtime_ipv6_multicast_enabled, runtime_ipv6_urpf_mode: .runtime_ipv6_urpf_mode, runtime_vrf: .runtime_vrf, runtime_ipv6_unicast_enabled: .runtime_ipv6_unicast_enabled, runtime_rmac_group: .runtime_rmac_group}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        l3_metadata$vrf <= runtime_vrf;
        qos_metadata$outer_dscp <= l3_metadata$lkp_ip_tc;
        ipv6_metadata$ipv6_unicast_enabled <= runtime_ipv6_unicast_enabled;
        ipv6_metadata$ipv6_urpf_mode <= runtime_ipv6_urpf_mode;
        l3_metadata$rmac_group <= runtime_rmac_group;
        l2_metadata$lkp_mac_sa <= ethernet$srcAddr;
        l2_metadata$lkp_mac_da <= ethernet$dstAddr;
        l3_metadata$lkp_ip_type <= 'h2;
        ipv6_metadata$lkp_ipv6_sa <= inner_ipv6$srcAddr;
        ipv6_metadata$lkp_ipv6_da <= inner_ipv6$dstAddr;
        l3_metadata$lkp_ip_version <= inner_ipv6$version;
        l3_metadata$lkp_ip_tc <= inner_ipv6$trafficClass;
        multicast_metadata$bd_mrpf_group <= runtime_mrpf_group;
        multicast_metadata$ipv6_multicast_enabled <= runtime_ipv6_multicast_enabled;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_tunnel_inner_ipv6_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateTunnelInnerIpv6RspT {pkt: pkt, l3_metadata$rmac_group: l3_metadata$rmac_group, qos_metadata$outer_dscp: qos_metadata$outer_dscp, multicast_metadata$bd_mrpf_group: multicast_metadata$bd_mrpf_group, l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, l3_metadata$vrf: l3_metadata$vrf, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, ipv6_metadata$ipv6_unicast_enabled: ipv6_metadata$ipv6_unicast_enabled, ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa, ipv6_metadata$ipv6_urpf_mode: ipv6_metadata$ipv6_urpf_mode, ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, multicast_metadata$ipv6_multicast_enabled: multicast_metadata$ipv6_multicast_enabled, l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version, l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_TUNNEL_INNER_NON_IP ======

interface TerminateTunnelInnerNonIp;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateTunnelInnerNonIp  (TerminateTunnelInnerNonIp);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) acl_metadata$bd_label <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$bd_stats_idx <- mkReg(0);
  Reg#(Bit#(2)) l3_metadata$lkp_ip_type <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule terminate_tunnel_inner_non_ip_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateTunnelInnerNonIpReqT {pkt: .pkt, inner_ethernet$etherType: .inner_ethernet$etherType, runtime_bd_label: .runtime_bd_label, runtime_bd: .runtime_bd, runtime_stats_idx: .runtime_stats_idx}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        ingress_metadata$bd <= runtime_bd;
        acl_metadata$bd_label <= runtime_bd_label;
        l2_metadata$bd_stats_idx <= runtime_stats_idx;
        l3_metadata$lkp_ip_type <= 'h0;
        l2_metadata$lkp_mac_type <= inner_ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_tunnel_inner_non_ip_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateTunnelInnerNonIpRspT {pkt: pkt, l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type, ingress_metadata$bd: ingress_metadata$bd, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type, acl_metadata$bd_label: acl_metadata$bd_label, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, l2_metadata$bd_stats_idx: l2_metadata$bd_stats_idx};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TERMINATE_VPLS ======

interface TerminateVpls;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTerminateVpls  (TerminateVpls);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) tunnel_metadata$tunnel_terminate <- mkReg(0);
  Reg#(Bit#(5)) tunnel_metadata$ingress_tunnel_type <- mkReg(0);
  Reg#(Bit#(16)) ingress_metadata$bd <- mkReg(0);
  Reg#(Bit#(16)) l2_metadata$lkp_mac_type <- mkReg(0);
  rule terminate_vpls_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TerminateVplsReqT {pkt: .pkt, inner_ethernet$etherType: .inner_ethernet$etherType, runtime_tunnel_type: .runtime_tunnel_type, runtime_bd: .runtime_bd}: begin
        tunnel_metadata$tunnel_terminate <= 'h1;
        tunnel_metadata$ingress_tunnel_type <= runtime_tunnel_type;
        ingress_metadata$bd <= runtime_bd;
        l2_metadata$lkp_mac_type <= inner_ethernet$etherType;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule terminate_vpls_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TerminateVplsRspT {pkt: pkt, tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type, ingress_metadata$bd: ingress_metadata$bd};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TUNNEL_LOOKUP_MISS ======

interface TunnelLookupMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkATunnelLookupMiss  (ATunnelLookupMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule tunnel_lookup_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TunnelLookupMissReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule tunnel_lookup_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TunnelLookupMissRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TUNNEL_MTU_CHECK ======

interface TunnelMtuCheck;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTunnelMtuCheck  (TunnelMtuCheck);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule tunnel_mtu_check_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TunnelMtuCheckReqT {pkt: .pkt, runtime_l3_mtu: .runtime_l3_mtu}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule tunnel_mtu_check_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TunnelMtuCheckRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== TUNNEL_MTU_MISS ======

interface TunnelMtuMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkTunnelMtuMiss  (TunnelMtuMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(16)) l3_metadata$l3_mtu_check <- mkReg(0);
  rule tunnel_mtu_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged TunnelMtuMissReqT {pkt: .pkt}: begin
        l3_metadata$l3_mtu_check <= 'hffff;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule tunnel_mtu_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged TunnelMtuMissRspT {pkt: pkt, l3_metadata$l3_mtu_check: l3_metadata$l3_mtu_check};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== UPDATE_INGRESS_BD_STATS ======

interface UpdateIngressBdStats;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkUpdateIngressBdStats  (UpdateIngressBdStats);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  rule update_ingress_bd_stats_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged UpdateIngressBdStatsReqT {pkt: .pkt}: begin
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule update_ingress_bd_stats_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged UpdateIngressBdStatsRspT {pkt: pkt};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== URPF_BD_MISS ======

interface UrpfBdMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkUrpfBdMiss  (UrpfBdMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$urpf_check_fail <- mkReg(0);
  rule urpf_bd_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged UrpfBdMissReqT {pkt: .pkt}: begin
        l3_metadata$urpf_check_fail <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule urpf_bd_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged UrpfBdMissRspT {pkt: pkt, l3_metadata$urpf_check_fail: l3_metadata$urpf_check_fail};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== URPF_MISS ======

interface UrpfMiss;
  interface Server#(BBRequest, BBResponse) prev_control_state;
endinterface
(* synthesize *)
module mkUrpfMiss  (UrpfMiss);
  RX #(BBRequest) rx_prev_control_state <- mkRX;
  TX #(BBResponse) tx_prev_control_state <- mkTX;
  let rx_info_prev_control_state = rx_prev_control_state.u;
  let tx_info_prev_control_state = tx_prev_control_state.u;
  FIFOF#(PacketInstance) curr_packet_ff <- mkFIFOF;
  Reg#(Bit#(1)) l3_metadata$urpf_check_fail <- mkReg(0);
  rule urpf_miss_request;
    let v = rx_info_prev_control_state.first;
    rx_info_prev_control_state.deq;
    case (v) matches
      tagged UrpfMissReqT {pkt: .pkt}: begin
        l3_metadata$urpf_check_fail <= 'h1;
        curr_packet_ff.enq(pkt);
      end
    endcase
  endrule

  rule urpf_miss_response;
    let pkt <- toGet(curr_packet_ff).get;
    BBResponse rsp = tagged UrpfMissRspT {pkt: pkt, l3_metadata$urpf_check_fail: l3_metadata$urpf_check_fail};
    tx_info_prev_control_state.enq(rsp);
  endrule

  interface prev_control_state = toServer(rx_prev_control_state.e, tx_prev_control_state.e);
endmodule

// ====== ACL_STATS ======

typedef struct {
} AclStatsReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_ACL_STATS,
  ACL_STATS_UPDATE
} AclStatsActionT deriving (Bits, Eq, FShow);
typedef struct {
  AclStatsActionT _action;
} AclStatsRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_acl_stats(Bit#(0) msgtype);
import "BDPI" function Action matchtable_write_acl_stats(Bit#(0) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(40, 0, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(40) id, Bit#(0) key);
    actionvalue
      let v <- matchtable_read_acl_stats(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(40) id, Bit#(0) key, Bit#(1) data);
    action
      matchtable_write_acl_stats(key, data);
    endaction
  endfunction

endinstance
interface AclStats;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkAclStats  (AclStats);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  FIFOF#(MetadataT) metadata_ff <- mkFIFOF;
  rule rl_handle_action_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    packet_ff.enq(pkt);
    metadata_ff.enq(meta);
    BBRequest req = tagged AclStatsUpdateReqT {pkt: pkt};
    bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
  endrule

  rule rl_handle_action_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff).get;
    case (v) matches
      tagged AclStatsUpdateRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged AclStatsAclStatsUpdateRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== BD_FLOOD ======

typedef struct {
  Bit#(8) padding;
  Bit#(16) ingress_metadata$bd;
  Bit#(3) l2_metadata$lkp_pkt_type;
} BdFloodReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_BD_FLOOD,
  NOP,
  SET_BD_FLOOD_MC_INDEX
} BdFloodActionT deriving (Bits, Eq, FShow);
typedef struct {
  BdFloodActionT _action;
  Bit#(16) runtime_mc_index;
} BdFloodRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_bd_flood(Bit#(27) msgtype);
import "BDPI" function Action matchtable_write_bd_flood(Bit#(27) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(55, 27, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(55) id, Bit#(27) key);
    actionvalue
      let v <- matchtable_read_bd_flood(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(55) id, Bit#(27) key, Bit#(18) data);
    action
      matchtable_write_bd_flood(key, data);
    endaction
  endfunction

endinstance
interface BdFlood;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkBdFlood  (BdFlood);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(55, 1024, SizeOf#(BdFloodReqT), SizeOf#(BdFloodRspT)) matchTable <- mkMatchTable("bd_flood.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    let l2_metadata$lkp_pkt_type = fromMaybe(?, meta.l2_metadata$lkp_pkt_type);
    BdFloodReqT req = BdFloodReqT {ingress_metadata$bd: ingress_metadata$bd,l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      BdFloodRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_BD_FLOOD_MC_INDEX: begin
          BBRequest req = tagged SetBdFloodMcIndexReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged BdFloodNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetBdFloodMcIndexRspT {pkt: .pkt, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged BdFloodSetBdFloodMcIndexRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== COMPUTE_IPV4_HASHES ======

typedef struct {
  Bit#(8) padding;
  Bit#(1) ingress_metadata$drop_flag;
} ComputeIpv4HashesReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_COMPUTE_IPV4_HASHES,
  COMPUTE_LKP_IPV4_HASH
} ComputeIpv4HashesActionT deriving (Bits, Eq, FShow);
typedef struct {
  ComputeIpv4HashesActionT _action;
} ComputeIpv4HashesRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_compute_ipv4_hashes(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_compute_ipv4_hashes(Bit#(9) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(70, 9, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(70) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_compute_ipv4_hashes(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(70) id, Bit#(9) key, Bit#(1) data);
    action
      matchtable_write_compute_ipv4_hashes(key, data);
    endaction
  endfunction

endinstance
interface ComputeIpv4Hashes;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkComputeIpv4Hashes  (ComputeIpv4Hashes);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(70, 256, SizeOf#(ComputeIpv4HashesReqT), SizeOf#(ComputeIpv4HashesRspT)) matchTable <- mkMatchTable("compute_ipv4_hashes.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
    ComputeIpv4HashesReqT req = ComputeIpv4HashesReqT {ingress_metadata$drop_flag: ingress_metadata$drop_flag};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ComputeIpv4HashesRspT resp = unpack(data);
      case (resp._action) matches
        COMPUTE_LKP_IPV4_HASH: begin
          BBRequest req = tagged ComputeLkpIpv4HashReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged ComputeLkpIpv4HashRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged ComputeIpv4HashesComputeLkpIpv4HashRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== COMPUTE_IPV6_HASHES ======

typedef struct {
  Bit#(8) padding;
  Bit#(1) ingress_metadata$drop_flag;
} ComputeIpv6HashesReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_COMPUTE_IPV6_HASHES,
  COMPUTE_LKP_IPV6_HASH
} ComputeIpv6HashesActionT deriving (Bits, Eq, FShow);
typedef struct {
  ComputeIpv6HashesActionT _action;
} ComputeIpv6HashesRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_compute_ipv6_hashes(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_compute_ipv6_hashes(Bit#(9) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(71, 9, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(71) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_compute_ipv6_hashes(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(71) id, Bit#(9) key, Bit#(1) data);
    action
      matchtable_write_compute_ipv6_hashes(key, data);
    endaction
  endfunction

endinstance
interface ComputeIpv6Hashes;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkComputeIpv6Hashes  (ComputeIpv6Hashes);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(71, 256, SizeOf#(ComputeIpv6HashesReqT), SizeOf#(ComputeIpv6HashesRspT)) matchTable <- mkMatchTable("compute_ipv6_hashes.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
    ComputeIpv6HashesReqT req = ComputeIpv6HashesReqT {ingress_metadata$drop_flag: ingress_metadata$drop_flag};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ComputeIpv6HashesRspT resp = unpack(data);
      case (resp._action) matches
        COMPUTE_LKP_IPV6_HASH: begin
          BBRequest req = tagged ComputeLkpIpv6HashReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged ComputeLkpIpv6HashRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged ComputeIpv6HashesComputeLkpIpv6HashRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== COMPUTE_NON_IP_HASHES ======

typedef struct {
  Bit#(8) padding;
  Bit#(1) ingress_metadata$drop_flag;
} ComputeNonIpHashesReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_COMPUTE_NON_IP_HASHES,
  COMPUTE_LKP_NON_IP_HASH
} ComputeNonIpHashesActionT deriving (Bits, Eq, FShow);
typedef struct {
  ComputeNonIpHashesActionT _action;
} ComputeNonIpHashesRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_compute_non_ip_hashes(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_compute_non_ip_hashes(Bit#(9) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(72, 9, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(72) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_compute_non_ip_hashes(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(72) id, Bit#(9) key, Bit#(1) data);
    action
      matchtable_write_compute_non_ip_hashes(key, data);
    endaction
  endfunction

endinstance
interface ComputeNonIpHashes;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkComputeNonIpHashes  (ComputeNonIpHashes);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(72, 256, SizeOf#(ComputeNonIpHashesReqT), SizeOf#(ComputeNonIpHashesRspT)) matchTable <- mkMatchTable("compute_non_ip_hashes.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
    ComputeNonIpHashesReqT req = ComputeNonIpHashesReqT {ingress_metadata$drop_flag: ingress_metadata$drop_flag};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ComputeNonIpHashesRspT resp = unpack(data);
      case (resp._action) matches
        COMPUTE_LKP_NON_IP_HASH: begin
          BBRequest req = tagged ComputeLkpNonIpHashReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged ComputeLkpNonIpHashRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged ComputeNonIpHashesComputeLkpNonIpHashRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== COMPUTE_OTHER_HASHES ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) hash_metadata$hash1;
} ComputeOtherHashesReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_COMPUTE_OTHER_HASHES,
  COMPUTED_TWO_HASHES,
  COMPUTED_ONE_HASH
} ComputeOtherHashesActionT deriving (Bits, Eq, FShow);
typedef struct {
  ComputeOtherHashesActionT _action;
} ComputeOtherHashesRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_compute_other_hashes(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_compute_other_hashes(Bit#(18) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(73, 18, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(73) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_compute_other_hashes(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(73) id, Bit#(18) key, Bit#(2) data);
    action
      matchtable_write_compute_other_hashes(key, data);
    endaction
  endfunction

endinstance
interface ComputeOtherHashes;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkComputeOtherHashes  (ComputeOtherHashes);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(73, 256, SizeOf#(ComputeOtherHashesReqT), SizeOf#(ComputeOtherHashesRspT)) matchTable <- mkMatchTable("compute_other_hashes.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let hash_metadata$hash1 = fromMaybe(?, meta.hash_metadata$hash1);
    ComputeOtherHashesReqT req = ComputeOtherHashesReqT {hash_metadata$hash1: hash_metadata$hash1};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ComputeOtherHashesRspT resp = unpack(data);
      case (resp._action) matches
        COMPUTED_TWO_HASHES: begin
          BBRequest req = tagged ComputedTwoHashesReqT {pkt: pkt, hash_metadata$hash1: hash_metadata$hash1, hash_metadata$hash2: hash_metadata$hash2};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        COMPUTED_ONE_HASH: begin
          BBRequest req = tagged ComputedOneHashReqT {pkt: pkt, hash_metadata$hash2: hash_metadata$hash2};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged ComputedTwoHashesRspT {pkt: .pkt, hash_metadata$entropy_hash: .hash_metadata$entropy_hash, intrinsic_metadata$mcast_hash: .intrinsic_metadata$mcast_hash}: begin
        meta.hash_metadata$entropy_hash = tagged Valid hash_metadata$entropy_hash;
        meta.intrinsic_metadata$mcast_hash = tagged Valid intrinsic_metadata$mcast_hash;
        MetadataResponse rsp = tagged ComputeOtherHashesComputedTwoHashesRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged ComputedOneHashRspT {pkt: .pkt, hash_metadata$entropy_hash: .hash_metadata$entropy_hash, intrinsic_metadata$mcast_hash: .intrinsic_metadata$mcast_hash, hash_metadata$hash1: .hash_metadata$hash1}: begin
        meta.hash_metadata$entropy_hash = tagged Valid hash_metadata$entropy_hash;
        meta.intrinsic_metadata$mcast_hash = tagged Valid intrinsic_metadata$mcast_hash;
        meta.hash_metadata$hash1 = tagged Valid hash_metadata$hash1;
        MetadataResponse rsp = tagged ComputeOtherHashesComputedOneHashRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== DMAC ======

typedef struct {
  Bit#(8) padding;
  Bit#(16) ingress_metadata$bd;
  Bit#(48) l2_metadata$lkp_mac_da;
} DmacReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_DMAC,
  NOP,
  DMAC_HIT,
  DMAC_MULTICAST_HIT,
  DMAC_MISS,
  DMAC_REDIRECT_NEXTHOP,
  DMAC_REDIRECT_ECMP,
  DMAC_DROP
} DmacActionT deriving (Bits, Eq, FShow);
typedef struct {
  DmacActionT _action;
  Bit#(16) runtime_ifindex;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} DmacRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(67)) matchtable_read_dmac(Bit#(72) msgtype);
import "BDPI" function Action matchtable_write_dmac(Bit#(72) msgtype, Bit#(67) data);
`endif
instance MatchTableSim#(9, 72, 67);
  function ActionValue#(Bit#(67)) matchtable_read(Bit#(9) id, Bit#(72) key);
    actionvalue
      let v <- matchtable_read_dmac(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(9) id, Bit#(72) key, Bit#(67) data);
    action
      matchtable_write_dmac(key, data);
    endaction
  endfunction

endinstance
interface Dmac;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
endinterface
(* synthesize *)
module mkDmac  (Dmac);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(7, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(7, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(9, 1024, SizeOf#(DmacReqT), SizeOf#(DmacRspT)) matchTable <- mkMatchTable("dmac.dat");
  Vector#(7, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(7) readyChannel = -1;
  for (Integer i=6; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    let l2_metadata$lkp_mac_da = fromMaybe(?, meta.l2_metadata$lkp_mac_da);
    DmacReqT req = DmacReqT {ingress_metadata$bd: ingress_metadata$bd,l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      DmacRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        DMAC_HIT: begin
          BBRequest req = tagged DmacHitReqT {pkt: pkt, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        DMAC_MULTICAST_HIT: begin
          BBRequest req = tagged DmacMulticastHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        DMAC_MISS: begin
          BBRequest req = tagged DmacMissReqT {pkt: pkt};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        DMAC_REDIRECT_NEXTHOP: begin
          BBRequest req = tagged DmacRedirectNexthopReqT {pkt: pkt, runtime_nexthop_index: resp.runtime_nexthop_index};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        DMAC_REDIRECT_ECMP: begin
          BBRequest req = tagged DmacRedirectEcmpReqT {pkt: pkt, runtime_ecmp_index: resp.runtime_ecmp_index};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        DMAC_DROP: begin
          BBRequest req = tagged DmacDropReqT {pkt: pkt};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged DmacNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DmacHitRspT {pkt: .pkt, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged DmacDmacHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DmacMulticastHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged DmacDmacMulticastHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DmacMissRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged DmacDmacMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DmacRedirectNexthopRspT {pkt: .pkt, l2_metadata$l2_redirect: .l2_metadata$l2_redirect, l2_metadata$l2_nexthop: .l2_metadata$l2_nexthop, l2_metadata$l2_nexthop_type: .l2_metadata$l2_nexthop_type}: begin
        meta.l2_metadata$l2_redirect = tagged Valid l2_metadata$l2_redirect;
        meta.l2_metadata$l2_nexthop = tagged Valid l2_metadata$l2_nexthop;
        meta.l2_metadata$l2_nexthop_type = tagged Valid l2_metadata$l2_nexthop_type;
        MetadataResponse rsp = tagged DmacDmacRedirectNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DmacRedirectEcmpRspT {pkt: .pkt, l2_metadata$l2_redirect: .l2_metadata$l2_redirect, l2_metadata$l2_nexthop: .l2_metadata$l2_nexthop, l2_metadata$l2_nexthop_type: .l2_metadata$l2_nexthop_type}: begin
        meta.l2_metadata$l2_redirect = tagged Valid l2_metadata$l2_redirect;
        meta.l2_metadata$l2_nexthop = tagged Valid l2_metadata$l2_nexthop;
        meta.l2_metadata$l2_nexthop_type = tagged Valid l2_metadata$l2_nexthop_type;
        MetadataResponse rsp = tagged DmacDmacRedirectEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DmacDropRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged DmacDmacDropRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
endmodule

// ====== DROP_STATS ======

typedef struct {
} DropStatsReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_DROP_STATS,
  DROP_STATS_UPDATE
} DropStatsActionT deriving (Bits, Eq, FShow);
typedef struct {
  DropStatsActionT _action;
} DropStatsRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_drop_stats(Bit#(0) msgtype);
import "BDPI" function Action matchtable_write_drop_stats(Bit#(0) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(42, 0, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(42) id, Bit#(0) key);
    actionvalue
      let v <- matchtable_read_drop_stats(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(42) id, Bit#(0) key, Bit#(1) data);
    action
      matchtable_write_drop_stats(key, data);
    endaction
  endfunction

endinstance
interface DropStats;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkDropStats  (DropStats);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  FIFOF#(MetadataT) metadata_ff <- mkFIFOF;
  rule rl_handle_action_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    packet_ff.enq(pkt);
    metadata_ff.enq(meta);
    BBRequest req = tagged DropStatsUpdateReqT {pkt: pkt};
    bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
  endrule

  rule rl_handle_action_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff).get;
    case (v) matches
      tagged DropStatsUpdateRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged DropStatsDropStatsUpdateRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== ECMP_GROUP ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) l3_metadata$nexthop_index;
} EcmpGroupReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_ECMP_GROUP,
  NOP,
  SET_ECMP_NEXTHOP_DETAILS,
  SET_ECMP_NEXTHOP_DETAILS_FOR_POST_ROUTED_FLOOD
} EcmpGroupActionT deriving (Bits, Eq, FShow);
typedef struct {
  EcmpGroupActionT _action;
  Bit#(16) runtime_ifindex;
  Bit#(16) runtime_bd;
  Bit#(16) runtime_nhop_index;
  Bit#(1) runtime_tunnel;
  Bit#(16) runtime_uuc_mc_index;
} EcmpGroupRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(67)) matchtable_read_ecmp_group(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_ecmp_group(Bit#(18) msgtype, Bit#(67) data);
`endif
instance MatchTableSim#(57, 18, 67);
  function ActionValue#(Bit#(67)) matchtable_read(Bit#(57) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_ecmp_group(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(57) id, Bit#(18) key, Bit#(67) data);
    action
      matchtable_write_ecmp_group(key, data);
    endaction
  endfunction

endinstance
interface EcmpGroup;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkEcmpGroup  (EcmpGroup);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(57, 1024, SizeOf#(EcmpGroupReqT), SizeOf#(EcmpGroupRspT)) matchTable <- mkMatchTable("ecmp_group.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
    EcmpGroupReqT req = EcmpGroupReqT {l3_metadata$nexthop_index: l3_metadata$nexthop_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      EcmpGroupRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_ECMP_NEXTHOP_DETAILS: begin
          BBRequest req = tagged SetEcmpNexthopDetailsReqT {pkt: pkt, runtime_bd: resp.runtime_bd, runtime_nhop_index: resp.runtime_nhop_index, runtime_ifindex: resp.runtime_ifindex, runtime_tunnel: resp.runtime_tunnel};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_ECMP_NEXTHOP_DETAILS_FOR_POST_ROUTED_FLOOD: begin
          BBRequest req = tagged SetEcmpNexthopDetailsForPostRoutedFloodReqT {pkt: pkt, runtime_uuc_mc_index: resp.runtime_uuc_mc_index, runtime_nhop_index: resp.runtime_nhop_index, runtime_bd: resp.runtime_bd};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged EcmpGroupNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetEcmpNexthopDetailsRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged EcmpGroupSetEcmpNexthopDetailsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetEcmpNexthopDetailsForPostRoutedFloodRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, fabric_metadata$dst_device: .fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged EcmpGroupSetEcmpNexthopDetailsForPostRoutedFloodRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== FABRIC_INGRESS_DST_LKP ======

typedef struct {
  Bit#(1) padding;
  Bit#(8) fabric_header$dstDevice;
} FabricIngressDstLkpReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_FABRIC_INGRESS_DST_LKP,
  NOP,
  TERMINATE_CPU_PACKET,
  SWITCH_FABRIC_UNICAST_PACKET,
  TERMINATE_FABRIC_UNICAST_PACKET,
  SWITCH_FABRIC_MULTICAST_PACKET,
  TERMINATE_FABRIC_MULTICAST_PACKET
} FabricIngressDstLkpActionT deriving (Bits, Eq, FShow);
typedef struct {
  FabricIngressDstLkpActionT _action;
} FabricIngressDstLkpRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(3)) matchtable_read_fabric_ingress_dst_lkp(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_fabric_ingress_dst_lkp(Bit#(9) msgtype, Bit#(3) data);
`endif
instance MatchTableSim#(63, 9, 3);
  function ActionValue#(Bit#(3)) matchtable_read(Bit#(63) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_fabric_ingress_dst_lkp(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(63) id, Bit#(9) key, Bit#(3) data);
    action
      matchtable_write_fabric_ingress_dst_lkp(key, data);
    endaction
  endfunction

endinstance
interface FabricIngressDstLkp;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
endinterface
(* synthesize *)
module mkFabricIngressDstLkp  (FabricIngressDstLkp);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(6, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(6, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(63, 256, SizeOf#(FabricIngressDstLkpReqT), SizeOf#(FabricIngressDstLkpRspT)) matchTable <- mkMatchTable("fabric_ingress_dst_lkp.dat");
  Vector#(6, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(6) readyChannel = -1;
  for (Integer i=5; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let fabric_header$dstDevice = fromMaybe(?, meta.fabric_header$dstDevice);
    FabricIngressDstLkpReqT req = FabricIngressDstLkpReqT {fabric_header$dstDevice: fabric_header$dstDevice};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      FabricIngressDstLkpRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_CPU_PACKET: begin
          BBRequest req = tagged TerminateCpuPacketReqT {pkt: pkt, fabric_payload_header$etherType: fabric_payload_header$etherType, fabric_header_cpu$txBypass: fabric_header_cpu$txBypass, fabric_header$dstPortOrGroup: fabric_header$dstPortOrGroup};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SWITCH_FABRIC_UNICAST_PACKET: begin
          BBRequest req = tagged SwitchFabricUnicastPacketReqT {pkt: pkt, fabric_header$dstDevice: fabric_header$dstDevice, fabric_header$dstPortOrGroup: fabric_header$dstPortOrGroup};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_FABRIC_UNICAST_PACKET: begin
          BBRequest req = tagged TerminateFabricUnicastPacketReqT {pkt: pkt, fabric_header_unicast$nexthopIndex: fabric_header_unicast$nexthopIndex, fabric_header_unicast$routed: fabric_header_unicast$routed, fabric_header_unicast$tunnelTerminate: fabric_header_unicast$tunnelTerminate, fabric_payload_header$etherType: fabric_payload_header$etherType, fabric_header_unicast$outerRouted: fabric_header_unicast$outerRouted, fabric_header_unicast$ingressTunnelType: fabric_header_unicast$ingressTunnelType, fabric_header$dstPortOrGroup: fabric_header$dstPortOrGroup};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        SWITCH_FABRIC_MULTICAST_PACKET: begin
          BBRequest req = tagged SwitchFabricMulticastPacketReqT {pkt: pkt, fabric_header$dstPortOrGroup: fabric_header$dstPortOrGroup};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_FABRIC_MULTICAST_PACKET: begin
          BBRequest req = tagged TerminateFabricMulticastPacketReqT {pkt: pkt, fabric_payload_header$etherType: fabric_payload_header$etherType, fabric_header_multicast$tunnelTerminate: fabric_header_multicast$tunnelTerminate, fabric_header_multicast$outerRouted: fabric_header_multicast$outerRouted, fabric_header_multicast$ingressTunnelType: fabric_header_multicast$ingressTunnelType, fabric_header_multicast$mcastGrp: fabric_header_multicast$mcastGrp, fabric_header_multicast$routed: fabric_header_multicast$routed};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged FabricIngressDstLkpNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateCpuPacketRspT {pkt: .pkt, egress_metadata$bypass: .egress_metadata$bypass, standard_metadata$egress_spec: .standard_metadata$egress_spec, ethernet$etherType: .ethernet$etherType}: begin
        meta.egress_metadata$bypass = tagged Valid egress_metadata$bypass;
        meta.standard_metadata$egress_spec = tagged Valid standard_metadata$egress_spec;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged FabricIngressDstLkpTerminateCpuPacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SwitchFabricUnicastPacketRspT {pkt: .pkt, fabric_metadata$fabric_header_present: .fabric_metadata$fabric_header_present, fabric_metadata$dst_port: .fabric_metadata$dst_port, fabric_metadata$dst_device: .fabric_metadata$dst_device}: begin
        meta.fabric_metadata$fabric_header_present = tagged Valid fabric_metadata$fabric_header_present;
        meta.fabric_metadata$dst_port = tagged Valid fabric_metadata$dst_port;
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        MetadataResponse rsp = tagged FabricIngressDstLkpSwitchFabricUnicastPacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateFabricUnicastPacketRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, tunnel_metadata$ingress_tunnel_type: .tunnel_metadata$ingress_tunnel_type, standard_metadata$egress_spec: .standard_metadata$egress_spec, l3_metadata$routed: .l3_metadata$routed, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, ethernet$etherType: .ethernet$etherType, l3_metadata$outer_routed: .l3_metadata$outer_routed}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        meta.tunnel_metadata$ingress_tunnel_type = tagged Valid tunnel_metadata$ingress_tunnel_type;
        meta.standard_metadata$egress_spec = tagged Valid standard_metadata$egress_spec;
        meta.l3_metadata$routed = tagged Valid l3_metadata$routed;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.l3_metadata$outer_routed = tagged Valid l3_metadata$outer_routed;
        MetadataResponse rsp = tagged FabricIngressDstLkpTerminateFabricUnicastPacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SwitchFabricMulticastPacketRspT {pkt: .pkt, fabric_metadata$fabric_header_present: .fabric_metadata$fabric_header_present, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$fabric_header_present = tagged Valid fabric_metadata$fabric_header_present;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged FabricIngressDstLkpSwitchFabricMulticastPacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateFabricMulticastPacketRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, tunnel_metadata$ingress_tunnel_type: .tunnel_metadata$ingress_tunnel_type, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l3_metadata$routed: .l3_metadata$routed, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, ethernet$etherType: .ethernet$etherType, l3_metadata$outer_routed: .l3_metadata$outer_routed}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        meta.tunnel_metadata$ingress_tunnel_type = tagged Valid tunnel_metadata$ingress_tunnel_type;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l3_metadata$routed = tagged Valid l3_metadata$routed;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.l3_metadata$outer_routed = tagged Valid l3_metadata$outer_routed;
        MetadataResponse rsp = tagged FabricIngressDstLkpTerminateFabricMulticastPacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
endmodule

// ====== FABRIC_INGRESS_SRC_LKP ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) fabric_header_multicast$ingressIfindex;
} FabricIngressSrcLkpReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_FABRIC_INGRESS_SRC_LKP,
  NOP,
  SET_INGRESS_IFINDEX_PROPERTIES
} FabricIngressSrcLkpActionT deriving (Bits, Eq, FShow);
typedef struct {
  FabricIngressSrcLkpActionT _action;
} FabricIngressSrcLkpRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_fabric_ingress_src_lkp(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_fabric_ingress_src_lkp(Bit#(18) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(64, 18, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(64) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_fabric_ingress_src_lkp(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(64) id, Bit#(18) key, Bit#(2) data);
    action
      matchtable_write_fabric_ingress_src_lkp(key, data);
    endaction
  endfunction

endinstance
interface FabricIngressSrcLkp;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkFabricIngressSrcLkp  (FabricIngressSrcLkp);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(64, 1024, SizeOf#(FabricIngressSrcLkpReqT), SizeOf#(FabricIngressSrcLkpRspT)) matchTable <- mkMatchTable("fabric_ingress_src_lkp.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let fabric_header_multicast$ingressIfindex = fromMaybe(?, meta.fabric_header_multicast$ingressIfindex);
    FabricIngressSrcLkpReqT req = FabricIngressSrcLkpReqT {fabric_header_multicast$ingressIfindex: fabric_header_multicast$ingressIfindex};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      FabricIngressSrcLkpRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_INGRESS_IFINDEX_PROPERTIES: begin
          BBRequest req = tagged SetIngressIfindexPropertiesReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged FabricIngressSrcLkpNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetIngressIfindexPropertiesRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged FabricIngressSrcLkpSetIngressIfindexPropertiesRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== FABRIC_LAG ======

typedef struct {
  Bit#(1) padding;
  Bit#(8) fabric_metadata$dst_device;
} FabricLagReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_FABRIC_LAG,
  NOP,
  SET_FABRIC_LAG_PORT,
  SET_FABRIC_MULTICAST
} FabricLagActionT deriving (Bits, Eq, FShow);
typedef struct {
  FabricLagActionT _action;
  Bit#(9) runtime_port;
} FabricLagRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(11)) matchtable_read_fabric_lag(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_fabric_lag(Bit#(9) msgtype, Bit#(11) data);
`endif
instance MatchTableSim#(66, 9, 11);
  function ActionValue#(Bit#(11)) matchtable_read(Bit#(66) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_fabric_lag(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(66) id, Bit#(9) key, Bit#(11) data);
    action
      matchtable_write_fabric_lag(key, data);
    endaction
  endfunction

endinstance
interface FabricLag;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkFabricLag  (FabricLag);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(66, 256, SizeOf#(FabricLagReqT), SizeOf#(FabricLagRspT)) matchTable <- mkMatchTable("fabric_lag.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let fabric_metadata$dst_device = fromMaybe(?, meta.fabric_metadata$dst_device);
    FabricLagReqT req = FabricLagReqT {fabric_metadata$dst_device: fabric_metadata$dst_device};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      FabricLagRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_FABRIC_LAG_PORT: begin
          BBRequest req = tagged SetFabricLagPortReqT {pkt: pkt, runtime_port: resp.runtime_port};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_FABRIC_MULTICAST: begin
          BBRequest req = tagged SetFabricMulticastReqT {pkt: pkt, intrinsic_metadata$mcast_grp: intrinsic_metadata$mcast_grp};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged FabricLagNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetFabricLagPortRspT {pkt: .pkt, standard_metadata$egress_spec: .standard_metadata$egress_spec}: begin
        meta.standard_metadata$egress_spec = tagged Valid standard_metadata$egress_spec;
        MetadataResponse rsp = tagged FabricLagSetFabricLagPortRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetFabricMulticastRspT {pkt: .pkt, multicast_metadata$mcast_grp: .multicast_metadata$mcast_grp}: begin
        meta.multicast_metadata$mcast_grp = tagged Valid multicast_metadata$mcast_grp;
        MetadataResponse rsp = tagged FabricLagSetFabricMulticastRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== FWD_RESULT ======

typedef struct {
  Bit#(4) padding;
  Bit#(1) l2_metadata$l2_redirect;
  Bit#(1) acl_metadata$acl_redirect;
  Bit#(1) acl_metadata$racl_redirect;
  Bit#(1) l3_metadata$rmac_hit;
  Bit#(1) l3_metadata$fib_hit;
  Bit#(3) l2_metadata$lkp_pkt_type;
  Bit#(2) l3_metadata$lkp_ip_type;
  Bit#(1) multicast_metadata$igmp_snooping_enabled;
  Bit#(1) multicast_metadata$mld_snooping_enabled;
  Bit#(1) multicast_metadata$mcast_route_hit;
  Bit#(1) multicast_metadata$mcast_bridge_hit;
  Bit#(16) multicast_metadata$mcast_rpf_group;
  Bit#(2) multicast_metadata$mcast_mode;
} FwdResultReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_FWD_RESULT,
  NOP,
  SET_L2_REDIRECT_ACTION,
  SET_FIB_REDIRECT_ACTION,
  SET_CPU_REDIRECT_ACTION,
  SET_ACL_REDIRECT_ACTION,
  SET_RACL_REDIRECT_ACTION,
  SET_MULTICAST_ROUTE_ACTION,
  SET_MULTICAST_BRIDGE_ACTION,
  SET_MULTICAST_FLOOD,
  SET_MULTICAST_DROP
} FwdResultActionT deriving (Bits, Eq, FShow);
typedef struct {
  FwdResultActionT _action;
} FwdResultRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(4)) matchtable_read_fwd_result(Bit#(36) msgtype);
import "BDPI" function Action matchtable_write_fwd_result(Bit#(36) msgtype, Bit#(4) data);
`endif
instance MatchTableSim#(56, 36, 4);
  function ActionValue#(Bit#(4)) matchtable_read(Bit#(56) id, Bit#(36) key);
    actionvalue
      let v <- matchtable_read_fwd_result(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(56) id, Bit#(36) key, Bit#(4) data);
    action
      matchtable_write_fwd_result(key, data);
    endaction
  endfunction

endinstance
interface FwdResult;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
  interface Client #(BBRequest, BBResponse) next_control_state_9;
endinterface
(* synthesize *)
module mkFwdResult  (FwdResult);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(10, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(10, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(56, 512, SizeOf#(FwdResultReqT), SizeOf#(FwdResultRspT)) matchTable <- mkMatchTable("fwd_result.dat");
  Vector#(10, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(10) readyChannel = -1;
  for (Integer i=9; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l2_metadata$l2_redirect = fromMaybe(?, meta.l2_metadata$l2_redirect);
    let acl_metadata$acl_redirect = fromMaybe(?, meta.acl_metadata$acl_redirect);
    let acl_metadata$racl_redirect = fromMaybe(?, meta.acl_metadata$racl_redirect);
    let l3_metadata$rmac_hit = fromMaybe(?, meta.l3_metadata$rmac_hit);
    let l3_metadata$fib_hit = fromMaybe(?, meta.l3_metadata$fib_hit);
    let l2_metadata$lkp_pkt_type = fromMaybe(?, meta.l2_metadata$lkp_pkt_type);
    let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
    let multicast_metadata$igmp_snooping_enabled = fromMaybe(?, meta.multicast_metadata$igmp_snooping_enabled);
    let multicast_metadata$mld_snooping_enabled = fromMaybe(?, meta.multicast_metadata$mld_snooping_enabled);
    let multicast_metadata$mcast_route_hit = fromMaybe(?, meta.multicast_metadata$mcast_route_hit);
    let multicast_metadata$mcast_bridge_hit = fromMaybe(?, meta.multicast_metadata$mcast_bridge_hit);
    let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
    let multicast_metadata$mcast_mode = fromMaybe(?, meta.multicast_metadata$mcast_mode);
    FwdResultReqT req = FwdResultReqT {l2_metadata$l2_redirect: l2_metadata$l2_redirect,acl_metadata$acl_redirect: acl_metadata$acl_redirect,acl_metadata$racl_redirect: acl_metadata$racl_redirect,l3_metadata$rmac_hit: l3_metadata$rmac_hit,l3_metadata$fib_hit: l3_metadata$fib_hit,l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type,l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type,multicast_metadata$igmp_snooping_enabled: multicast_metadata$igmp_snooping_enabled,multicast_metadata$mld_snooping_enabled: multicast_metadata$mld_snooping_enabled,multicast_metadata$mcast_route_hit: multicast_metadata$mcast_route_hit,multicast_metadata$mcast_bridge_hit: multicast_metadata$mcast_bridge_hit,multicast_metadata$mcast_rpf_group: multicast_metadata$mcast_rpf_group,multicast_metadata$mcast_mode: multicast_metadata$mcast_mode};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      FwdResultRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_L2_REDIRECT_ACTION: begin
          BBRequest req = tagged SetL2RedirectActionReqT {pkt: pkt, l2_metadata$l2_nexthop: l2_metadata$l2_nexthop, l2_metadata$l2_nexthop_type: l2_metadata$l2_nexthop_type};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_FIB_REDIRECT_ACTION: begin
          BBRequest req = tagged SetFibRedirectActionReqT {pkt: pkt, l3_metadata$fib_nexthop: l3_metadata$fib_nexthop, l3_metadata$fib_nexthop_type: l3_metadata$fib_nexthop_type};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        SET_CPU_REDIRECT_ACTION: begin
          BBRequest req = tagged SetCpuRedirectActionReqT {pkt: pkt};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        SET_ACL_REDIRECT_ACTION: begin
          BBRequest req = tagged SetAclRedirectActionReqT {pkt: pkt, acl_metadata$acl_nexthop: acl_metadata$acl_nexthop, acl_metadata$acl_nexthop_type: acl_metadata$acl_nexthop_type};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        SET_RACL_REDIRECT_ACTION: begin
          BBRequest req = tagged SetRaclRedirectActionReqT {pkt: pkt, acl_metadata$racl_nexthop: acl_metadata$racl_nexthop, acl_metadata$racl_nexthop_type: acl_metadata$racl_nexthop_type};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        SET_MULTICAST_ROUTE_ACTION: begin
          BBRequest req = tagged SetMulticastRouteActionReqT {pkt: pkt, multicast_metadata$multicast_route_mc_index: multicast_metadata$multicast_route_mc_index};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        SET_MULTICAST_BRIDGE_ACTION: begin
          BBRequest req = tagged SetMulticastBridgeActionReqT {pkt: pkt, multicast_metadata$multicast_bridge_mc_index: multicast_metadata$multicast_bridge_mc_index};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        SET_MULTICAST_FLOOD: begin
          BBRequest req = tagged SetMulticastFloodReqT {pkt: pkt};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
        SET_MULTICAST_DROP: begin
          BBRequest req = tagged SetMulticastDropReqT {pkt: pkt};
          bbReqFifo[9].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged FwdResultNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetL2RedirectActionRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, nexthop_metadata$nexthop_type: .nexthop_metadata$nexthop_type, fabric_metadata$dst_device: .fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        meta.nexthop_metadata$nexthop_type = tagged Valid nexthop_metadata$nexthop_type;
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged FwdResultSetL2RedirectActionRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetFibRedirectActionRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, nexthop_metadata$nexthop_type: .nexthop_metadata$nexthop_type, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l3_metadata$routed: .l3_metadata$routed, fabric_metadata$dst_device: .fabric_metadata$dst_device, fabric_metadata$reason_code: .fabric_metadata$reason_code}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        meta.nexthop_metadata$nexthop_type = tagged Valid nexthop_metadata$nexthop_type;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l3_metadata$routed = tagged Valid l3_metadata$routed;
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        MetadataResponse rsp = tagged FwdResultSetFibRedirectActionRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetCpuRedirectActionRspT {pkt: .pkt, l3_metadata$routed: .l3_metadata$routed, fabric_metadata$dst_device: .fabric_metadata$dst_device, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, standard_metadata$egress_spec: .standard_metadata$egress_spec}: begin
        meta.l3_metadata$routed = tagged Valid l3_metadata$routed;
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.standard_metadata$egress_spec = tagged Valid standard_metadata$egress_spec;
        MetadataResponse rsp = tagged FwdResultSetCpuRedirectActionRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetAclRedirectActionRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, nexthop_metadata$nexthop_type: .nexthop_metadata$nexthop_type, fabric_metadata$dst_device: .fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        meta.nexthop_metadata$nexthop_type = tagged Valid nexthop_metadata$nexthop_type;
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged FwdResultSetAclRedirectActionRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetRaclRedirectActionRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index, nexthop_metadata$nexthop_type: .nexthop_metadata$nexthop_type, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex, l3_metadata$routed: .l3_metadata$routed, fabric_metadata$dst_device: .fabric_metadata$dst_device}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        meta.nexthop_metadata$nexthop_type = tagged Valid nexthop_metadata$nexthop_type;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        meta.l3_metadata$routed = tagged Valid l3_metadata$routed;
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        MetadataResponse rsp = tagged FwdResultSetRaclRedirectActionRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMulticastRouteActionRspT {pkt: .pkt, l3_metadata$routed: .l3_metadata$routed, fabric_metadata$dst_device: .fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l3_metadata$same_bd_check: .l3_metadata$same_bd_check, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.l3_metadata$routed = tagged Valid l3_metadata$routed;
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l3_metadata$same_bd_check = tagged Valid l3_metadata$same_bd_check;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged FwdResultSetMulticastRouteActionRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMulticastBridgeActionRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged FwdResultSetMulticastBridgeActionRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMulticastFloodRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged FwdResultSetMulticastFloodRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMulticastDropRspT {pkt: .pkt, ingress_metadata$drop_reason: .ingress_metadata$drop_reason, ingress_metadata$drop_flag: .ingress_metadata$drop_flag}: begin
        meta.ingress_metadata$drop_reason = tagged Valid ingress_metadata$drop_reason;
        meta.ingress_metadata$drop_flag = tagged Valid ingress_metadata$drop_flag;
        MetadataResponse rsp = tagged FwdResultSetMulticastDropRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
  interface next_control_state_9 = toClient(bbReqFifo[9], bbRspFifo[9]);
endmodule

// ====== INGRESS_BD_STATS ======

typedef struct {
} IngressBdStatsReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INGRESS_BD_STATS,
  UPDATE_INGRESS_BD_STATS
} IngressBdStatsActionT deriving (Bits, Eq, FShow);
typedef struct {
  IngressBdStatsActionT _action;
} IngressBdStatsRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_ingress_bd_stats(Bit#(0) msgtype);
import "BDPI" function Action matchtable_write_ingress_bd_stats(Bit#(0) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(5, 0, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(5) id, Bit#(0) key);
    actionvalue
      let v <- matchtable_read_ingress_bd_stats(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(5) id, Bit#(0) key, Bit#(1) data);
    action
      matchtable_write_ingress_bd_stats(key, data);
    endaction
  endfunction

endinstance
interface IngressBdStats;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkIngressBdStats  (IngressBdStats);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  FIFOF#(MetadataT) metadata_ff <- mkFIFOF;
  rule rl_handle_action_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    packet_ff.enq(pkt);
    metadata_ff.enq(meta);
    BBRequest req = tagged UpdateIngressBdStatsReqT {pkt: pkt};
    bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
  endrule

  rule rl_handle_action_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff).get;
    case (v) matches
      tagged UpdateIngressBdStatsRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IngressBdStatsUpdateIngressBdStatsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== INGRESS_PORT_MAPPING ======

typedef struct {
  Bit#(9) standard_metadata$ingress_port;
} IngressPortMappingReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INGRESS_PORT_MAPPING,
  SET_IFINDEX
} IngressPortMappingActionT deriving (Bits, Eq, FShow);
typedef struct {
  IngressPortMappingActionT _action;
  Bit#(16) runtime_ifindex;
  Bit#(2) runtime_port_type;
} IngressPortMappingRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(19)) matchtable_read_ingress_port_mapping(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_ingress_port_mapping(Bit#(9) msgtype, Bit#(19) data);
`endif
instance MatchTableSim#(2, 9, 19);
  function ActionValue#(Bit#(19)) matchtable_read(Bit#(2) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_ingress_port_mapping(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(2) id, Bit#(9) key, Bit#(19) data);
    action
      matchtable_write_ingress_port_mapping(key, data);
    endaction
  endfunction

endinstance
interface IngressPortMapping;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkIngressPortMapping  (IngressPortMapping);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(2, 512, SizeOf#(IngressPortMappingReqT), SizeOf#(IngressPortMappingRspT)) matchTable <- mkMatchTable("ingress_port_mapping.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let standard_metadata$ingress_port = fromMaybe(?, meta.standard_metadata$ingress_port);
    IngressPortMappingReqT req = IngressPortMappingReqT {standard_metadata$ingress_port: standard_metadata$ingress_port};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IngressPortMappingRspT resp = unpack(data);
      case (resp._action) matches
        SET_IFINDEX: begin
          BBRequest req = tagged SetIfindexReqT {pkt: pkt, runtime_port_type: resp.runtime_port_type, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetIfindexRspT {pkt: .pkt, ingress_metadata$port_type: .ingress_metadata$port_type, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        meta.ingress_metadata$port_type = tagged Valid ingress_metadata$port_type;
        meta.ingress_metadata$ifindex = tagged Valid ingress_metadata$ifindex;
        MetadataResponse rsp = tagged IngressPortMappingSetIfindexRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== INGRESS_PORT_PROPERTIES ======

typedef struct {
  Bit#(9) standard_metadata$ingress_port;
} IngressPortPropertiesReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INGRESS_PORT_PROPERTIES,
  SET_INGRESS_PORT_PROPERTIES
} IngressPortPropertiesActionT deriving (Bits, Eq, FShow);
typedef struct {
  IngressPortPropertiesActionT _action;
  Bit#(16) runtime_if_label;
} IngressPortPropertiesRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(17)) matchtable_read_ingress_port_properties(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_ingress_port_properties(Bit#(9) msgtype, Bit#(17) data);
`endif
instance MatchTableSim#(3, 9, 17);
  function ActionValue#(Bit#(17)) matchtable_read(Bit#(3) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_ingress_port_properties(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(3) id, Bit#(9) key, Bit#(17) data);
    action
      matchtable_write_ingress_port_properties(key, data);
    endaction
  endfunction

endinstance
interface IngressPortProperties;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkIngressPortProperties  (IngressPortProperties);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(3, 512, SizeOf#(IngressPortPropertiesReqT), SizeOf#(IngressPortPropertiesRspT)) matchTable <- mkMatchTable("ingress_port_properties.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let standard_metadata$ingress_port = fromMaybe(?, meta.standard_metadata$ingress_port);
    IngressPortPropertiesReqT req = IngressPortPropertiesReqT {standard_metadata$ingress_port: standard_metadata$ingress_port};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IngressPortPropertiesRspT resp = unpack(data);
      case (resp._action) matches
        SET_INGRESS_PORT_PROPERTIES: begin
          BBRequest req = tagged SetIngressPortPropertiesReqT {pkt: pkt, runtime_if_label: resp.runtime_if_label};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetIngressPortPropertiesRspT {pkt: .pkt, acl_metadata$if_label: .acl_metadata$if_label}: begin
        meta.acl_metadata$if_label = tagged Valid acl_metadata$if_label;
        MetadataResponse rsp = tagged IngressPortPropertiesSetIngressPortPropertiesRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== INT_SINK_UPDATE_OUTER ======

typedef struct {
  Bit#(6) padding;
  Bit#(Bool) valid_vxlan_gpe_int_header;
  Bit#(Bool) valid_ipv4;
  Bit#(1) int_metadata_i2e$sink;
} IntSinkUpdateOuterReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_SINK_UPDATE_OUTER,
  INT_SINK_UPDATE_VXLAN_GPE_V4,
  NOP
} IntSinkUpdateOuterActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntSinkUpdateOuterActionT _action;
} IntSinkUpdateOuterRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_int_sink_update_outer(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_int_sink_update_outer(Bit#(9) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(69, 9, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(69) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_int_sink_update_outer(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(69) id, Bit#(9) key, Bit#(2) data);
    action
      matchtable_write_int_sink_update_outer(key, data);
    endaction
  endfunction

endinstance
interface IntSinkUpdateOuter;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIntSinkUpdateOuter  (IntSinkUpdateOuter);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(69, 256, SizeOf#(IntSinkUpdateOuterReqT), SizeOf#(IntSinkUpdateOuterRspT)) matchTable <- mkMatchTable("int_sink_update_outer.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let v$x$l$a$n$_$g$p$e$_$i$n$t$_$h$e$a$d$e$r = fromMaybe(?, meta.v$x$l$a$n$_$g$p$e$_$i$n$t$_$h$e$a$d$e$r);
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let int_metadata_i2e$sink = fromMaybe(?, meta.int_metadata_i2e$sink);
    IntSinkUpdateOuterReqT req = IntSinkUpdateOuterReqT {v$x$l$a$n$_$g$p$e$_$i$n$t$_$h$e$a$d$e$r: v$x$l$a$n$_$g$p$e$_$i$n$t$_$h$e$a$d$e$r,i$p$v$4: i$p$v$4,int_metadata_i2e$sink: int_metadata_i2e$sink};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntSinkUpdateOuterRspT resp = unpack(data);
      case (resp._action) matches
        INT_SINK_UPDATE_VXLAN_GPE_V4: begin
          BBRequest req = tagged IntSinkUpdateVxlanGpeV4ReqT {pkt: pkt, vxlan_gpe_int_header$next_proto: vxlan_gpe_int_header$next_proto};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntSinkUpdateVxlanGpeV4RspT {pkt: .pkt, vxlan_gpe$next_proto: .vxlan_gpe$next_proto}: begin
        meta.vxlan_gpe$next_proto = tagged Valid vxlan_gpe$next_proto;
        MetadataResponse rsp = tagged IntSinkUpdateOuterIntSinkUpdateVxlanGpeV4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IntSinkUpdateOuterNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== INT_SOURCE ======

typedef struct {
  Bit#(4) padding;
  Bit#(Bool) valid_int_header;
  Bit#(Bool) valid_ipv4;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
  Bit#(Bool) valid_inner_ipv4;
  Bit#(32) inner_ipv4$dstAddr;
  Bit#(32) inner_ipv4$srcAddr;
} IntSourceReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_SOURCE,
  INT_SET_SRC,
  INT_SET_NO_SRC
} IntSourceActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntSourceActionT _action;
} IntSourceRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_int_source(Bit#(135) msgtype);
import "BDPI" function Action matchtable_write_int_source(Bit#(135) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(67, 135, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(67) id, Bit#(135) key);
    actionvalue
      let v <- matchtable_read_int_source(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(67) id, Bit#(135) key, Bit#(2) data);
    action
      matchtable_write_int_source(key, data);
    endaction
  endfunction

endinstance
interface IntSource;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIntSource  (IntSource);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(67, 256, SizeOf#(IntSourceReqT), SizeOf#(IntSourceRspT)) matchTable <- mkMatchTable("int_source.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$n$t$_$h$e$a$d$e$r = fromMaybe(?, meta.i$n$t$_$h$e$a$d$e$r);
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    let i$n$n$e$r$_$i$p$v$4 = fromMaybe(?, meta.i$n$n$e$r$_$i$p$v$4);
    let inner_ipv4$dstAddr = fromMaybe(?, meta.inner_ipv4$dstAddr);
    let inner_ipv4$srcAddr = fromMaybe(?, meta.inner_ipv4$srcAddr);
    IntSourceReqT req = IntSourceReqT {i$n$t$_$h$e$a$d$e$r: i$n$t$_$h$e$a$d$e$r,i$p$v$4: i$p$v$4,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa,i$n$n$e$r$_$i$p$v$4: i$n$n$e$r$_$i$p$v$4,inner_ipv4$dstAddr: inner_ipv4$dstAddr,inner_ipv4$srcAddr: inner_ipv4$srcAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntSourceRspT resp = unpack(data);
      case (resp._action) matches
        INT_SET_SRC: begin
          BBRequest req = tagged IntSetSrcReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_NO_SRC: begin
          BBRequest req = tagged IntSetNoSrcReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntSetSrcRspT {pkt: .pkt, int_metadata_i2e$source: .int_metadata_i2e$source}: begin
        meta.int_metadata_i2e$source = tagged Valid int_metadata_i2e$source;
        MetadataResponse rsp = tagged IntSourceIntSetSrcRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetNoSrcRspT {pkt: .pkt, int_metadata_i2e$source: .int_metadata_i2e$source}: begin
        meta.int_metadata_i2e$source = tagged Valid int_metadata_i2e$source;
        MetadataResponse rsp = tagged IntSourceIntSetNoSrcRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== INT_TERMINATE ======

typedef struct {
  Bit#(4) padding;
  Bit#(Bool) valid_int_header;
  Bit#(Bool) valid_vxlan_gpe_int_header;
  Bit#(Bool) valid_ipv4;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
  Bit#(Bool) valid_inner_ipv4;
  Bit#(32) inner_ipv4$dstAddr;
} IntTerminateReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_TERMINATE,
  INT_SINK_GPE,
  INT_NO_SINK
} IntTerminateActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntTerminateActionT _action;
  Bit#(32) runtime_mirror_id;
} IntTerminateRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_int_terminate(Bit#(72) msgtype);
import "BDPI" function Action matchtable_write_int_terminate(Bit#(72) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(68, 72, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(68) id, Bit#(72) key);
    actionvalue
      let v <- matchtable_read_int_terminate(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(68) id, Bit#(72) key, Bit#(34) data);
    action
      matchtable_write_int_terminate(key, data);
    endaction
  endfunction

endinstance
interface IntTerminate;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIntTerminate  (IntTerminate);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(68, 256, SizeOf#(IntTerminateReqT), SizeOf#(IntTerminateRspT)) matchTable <- mkMatchTable("int_terminate.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$n$t$_$h$e$a$d$e$r = fromMaybe(?, meta.i$n$t$_$h$e$a$d$e$r);
    let v$x$l$a$n$_$g$p$e$_$i$n$t$_$h$e$a$d$e$r = fromMaybe(?, meta.v$x$l$a$n$_$g$p$e$_$i$n$t$_$h$e$a$d$e$r);
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    let i$n$n$e$r$_$i$p$v$4 = fromMaybe(?, meta.i$n$n$e$r$_$i$p$v$4);
    let inner_ipv4$dstAddr = fromMaybe(?, meta.inner_ipv4$dstAddr);
    IntTerminateReqT req = IntTerminateReqT {i$n$t$_$h$e$a$d$e$r: i$n$t$_$h$e$a$d$e$r,v$x$l$a$n$_$g$p$e$_$i$n$t$_$h$e$a$d$e$r: v$x$l$a$n$_$g$p$e$_$i$n$t$_$h$e$a$d$e$r,i$p$v$4: i$p$v$4,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da,i$n$n$e$r$_$i$p$v$4: i$n$n$e$r$_$i$p$v$4,inner_ipv4$dstAddr: inner_ipv4$dstAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntTerminateRspT resp = unpack(data);
      case (resp._action) matches
        INT_SINK_GPE: begin
          BBRequest req = tagged IntSinkGpeReqT {pkt: pkt, runtime_mirror_id: resp.runtime_mirror_id};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INT_NO_SINK: begin
          BBRequest req = tagged IntNoSinkReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntSinkGpeRspT {pkt: .pkt, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id, int_metadata_i2e$sink: .int_metadata_i2e$sink}: begin
        meta.i2e_metadata$mirror_session_id = tagged Valid i2e_metadata$mirror_session_id;
        meta.int_metadata_i2e$sink = tagged Valid int_metadata_i2e$sink;
        MetadataResponse rsp = tagged IntTerminateIntSinkGpeRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntNoSinkRspT {pkt: .pkt, int_metadata_i2e$sink: .int_metadata_i2e$sink}: begin
        meta.int_metadata_i2e$sink = tagged Valid int_metadata_i2e$sink;
        MetadataResponse rsp = tagged IntTerminateIntNoSinkRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IP_ACL ======

typedef struct {
  Bit#(1) padding;
  Bit#(16) acl_metadata$if_label;
  Bit#(16) acl_metadata$bd_label;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
  Bit#(8) l3_metadata$lkp_ip_proto;
  Bit#(16) l3_metadata$lkp_l4_sport;
  Bit#(16) l3_metadata$lkp_l4_dport;
  Bit#(8) tcp$flags;
  Bit#(8) l3_metadata$lkp_ip_ttl;
} IpAclReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IP_ACL,
  NOP,
  ACL_DENY,
  ACL_PERMIT,
  ACL_MIRROR,
  ACL_REDIRECT_NEXTHOP,
  ACL_REDIRECT_ECMP
} IpAclActionT deriving (Bits, Eq, FShow);
typedef struct {
  IpAclActionT _action;
  Bit#(14) runtime_acl_stats_index;
  Bit#(16) runtime_acl_meter_index;
  Bit#(1) runtime_acl_copy;
  Bit#(16) runtime_acl_copy_reason;
  Bit#(32) runtime_session_id;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} IpAclRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(114)) matchtable_read_ip_acl(Bit#(153) msgtype);
import "BDPI" function Action matchtable_write_ip_acl(Bit#(153) msgtype, Bit#(114) data);
`endif
instance MatchTableSim#(35, 153, 114);
  function ActionValue#(Bit#(114)) matchtable_read(Bit#(35) id, Bit#(153) key);
    actionvalue
      let v <- matchtable_read_ip_acl(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(35) id, Bit#(153) key, Bit#(114) data);
    action
      matchtable_write_ip_acl(key, data);
    endaction
  endfunction

endinstance
interface IpAcl;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
endinterface
(* synthesize *)
module mkIpAcl  (IpAcl);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(6, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(6, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(35, 512, SizeOf#(IpAclReqT), SizeOf#(IpAclRspT)) matchTable <- mkMatchTable("ip_acl.dat");
  Vector#(6, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(6) readyChannel = -1;
  for (Integer i=5; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let acl_metadata$if_label = fromMaybe(?, meta.acl_metadata$if_label);
    let acl_metadata$bd_label = fromMaybe(?, meta.acl_metadata$bd_label);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    let l3_metadata$lkp_ip_proto = fromMaybe(?, meta.l3_metadata$lkp_ip_proto);
    let l3_metadata$lkp_l4_sport = fromMaybe(?, meta.l3_metadata$lkp_l4_sport);
    let l3_metadata$lkp_l4_dport = fromMaybe(?, meta.l3_metadata$lkp_l4_dport);
    let tcp$flags = fromMaybe(?, meta.tcp$flags);
    let l3_metadata$lkp_ip_ttl = fromMaybe(?, meta.l3_metadata$lkp_ip_ttl);
    IpAclReqT req = IpAclReqT {acl_metadata$if_label: acl_metadata$if_label,acl_metadata$bd_label: acl_metadata$bd_label,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da,l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto,l3_metadata$lkp_l4_sport: l3_metadata$lkp_l4_sport,l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport,tcp$flags: tcp$flags,l3_metadata$lkp_ip_ttl: l3_metadata$lkp_ip_ttl};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IpAclRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        ACL_DENY: begin
          BBRequest req = tagged AclDenyReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        ACL_PERMIT: begin
          BBRequest req = tagged AclPermitReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        ACL_MIRROR: begin
          BBRequest req = tagged AclMirrorReqT {pkt: pkt, intrinsic_metadata$ingress_global_tstamp: intrinsic_metadata$ingress_global_tstamp, runtime_session_id: resp.runtime_session_id, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        ACL_REDIRECT_NEXTHOP: begin
          BBRequest req = tagged AclRedirectNexthopReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_copy: resp.runtime_acl_copy, runtime_nexthop_index: resp.runtime_nexthop_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        ACL_REDIRECT_ECMP: begin
          BBRequest req = tagged AclRedirectEcmpReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_copy: resp.runtime_acl_copy, runtime_ecmp_index: resp.runtime_ecmp_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IpAclNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclDenyRspT {pkt: .pkt, acl_metadata$acl_deny: .acl_metadata$acl_deny, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_copy: .acl_metadata$acl_copy}: begin
        meta.acl_metadata$acl_deny = tagged Valid acl_metadata$acl_deny;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        MetadataResponse rsp = tagged IpAclAclDenyRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclPermitRspT {pkt: .pkt, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_copy: .acl_metadata$acl_copy}: begin
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        MetadataResponse rsp = tagged IpAclAclPermitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclMirrorRspT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id}: begin
        meta.i2e_metadata$ingress_tstamp = tagged Valid i2e_metadata$ingress_tstamp;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.i2e_metadata$mirror_session_id = tagged Valid i2e_metadata$mirror_session_id;
        MetadataResponse rsp = tagged IpAclAclMirrorRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclRedirectNexthopRspT {pkt: .pkt, meter_metadata$meter_index: .meter_metadata$meter_index, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$acl_redirect: .acl_metadata$acl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_nexthop: .acl_metadata$acl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_nexthop_type: .acl_metadata$acl_nexthop_type}: begin
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$acl_redirect = tagged Valid acl_metadata$acl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_nexthop = tagged Valid acl_metadata$acl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_nexthop_type = tagged Valid acl_metadata$acl_nexthop_type;
        MetadataResponse rsp = tagged IpAclAclRedirectNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclRedirectEcmpRspT {pkt: .pkt, meter_metadata$meter_index: .meter_metadata$meter_index, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$acl_redirect: .acl_metadata$acl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_nexthop: .acl_metadata$acl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_nexthop_type: .acl_metadata$acl_nexthop_type}: begin
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$acl_redirect = tagged Valid acl_metadata$acl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_nexthop = tagged Valid acl_metadata$acl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_nexthop_type = tagged Valid acl_metadata$acl_nexthop_type;
        MetadataResponse rsp = tagged IpAclAclRedirectEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
endmodule

// ====== IPSG ======

typedef struct {
  Bit#(5) padding;
  Bit#(16) ingress_metadata$ifindex;
  Bit#(16) ingress_metadata$bd;
  Bit#(48) l2_metadata$lkp_mac_sa;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
} IpsgReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPSG,
  ON_MISS
} IpsgActionT deriving (Bits, Eq, FShow);
typedef struct {
  IpsgActionT _action;
} IpsgRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_ipsg(Bit#(117) msgtype);
import "BDPI" function Action matchtable_write_ipsg(Bit#(117) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(62, 117, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(62) id, Bit#(117) key);
    actionvalue
      let v <- matchtable_read_ipsg(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(62) id, Bit#(117) key, Bit#(1) data);
    action
      matchtable_write_ipsg(key, data);
    endaction
  endfunction

endinstance
interface Ipsg;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkIpsg  (Ipsg);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(62, 1024, SizeOf#(IpsgReqT), SizeOf#(IpsgRspT)) matchTable <- mkMatchTable("ipsg.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$ifindex = fromMaybe(?, meta.ingress_metadata$ifindex);
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    let l2_metadata$lkp_mac_sa = fromMaybe(?, meta.l2_metadata$lkp_mac_sa);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    IpsgReqT req = IpsgReqT {ingress_metadata$ifindex: ingress_metadata$ifindex,ingress_metadata$bd: ingress_metadata$bd,l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IpsgRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IpsgOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== IPSG_PERMIT_SPECIAL ======

typedef struct {
  Bit#(7) padding;
  Bit#(8) l3_metadata$lkp_ip_proto;
  Bit#(16) l3_metadata$lkp_l4_dport;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
} IpsgPermitSpecialReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPSG_PERMIT_SPECIAL,
  IPSG_MISS
} IpsgPermitSpecialActionT deriving (Bits, Eq, FShow);
typedef struct {
  IpsgPermitSpecialActionT _action;
} IpsgPermitSpecialRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_ipsg_permit_special(Bit#(63) msgtype);
import "BDPI" function Action matchtable_write_ipsg_permit_special(Bit#(63) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(61, 63, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(61) id, Bit#(63) key);
    actionvalue
      let v <- matchtable_read_ipsg_permit_special(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(61) id, Bit#(63) key, Bit#(1) data);
    action
      matchtable_write_ipsg_permit_special(key, data);
    endaction
  endfunction

endinstance
interface IpsgPermitSpecial;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkIpsgPermitSpecial  (IpsgPermitSpecial);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(61, 512, SizeOf#(IpsgPermitSpecialReqT), SizeOf#(IpsgPermitSpecialRspT)) matchTable <- mkMatchTable("ipsg_permit_special.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$lkp_ip_proto = fromMaybe(?, meta.l3_metadata$lkp_ip_proto);
    let l3_metadata$lkp_l4_dport = fromMaybe(?, meta.l3_metadata$lkp_l4_dport);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    IpsgPermitSpecialReqT req = IpsgPermitSpecialReqT {l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto,l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IpsgPermitSpecialRspT resp = unpack(data);
      case (resp._action) matches
        IPSG_MISS: begin
          BBRequest req = tagged IpsgMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IpsgMissRspT {pkt: .pkt, security_metadata$ipsg_check_fail: .security_metadata$ipsg_check_fail}: begin
        meta.security_metadata$ipsg_check_fail = tagged Valid security_metadata$ipsg_check_fail;
        MetadataResponse rsp = tagged IpsgPermitSpecialIpsgMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== IPV4_DEST_VTEP ======

typedef struct {
  Bit#(1) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(32) ipv4$dstAddr;
  Bit#(5) tunnel_metadata$ingress_tunnel_type;
} Ipv4DestVtepReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_DEST_VTEP,
  NOP,
  SET_TUNNEL_TERMINATION_FLAG,
  SET_TUNNEL_VNI_AND_TERMINATION_FLAG
} Ipv4DestVtepActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4DestVtepActionT _action;
  Bit#(24) runtime_tunnel_vni;
} Ipv4DestVtepRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(26)) matchtable_read_ipv4_dest_vtep(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_ipv4_dest_vtep(Bit#(54) msgtype, Bit#(26) data);
`endif
instance MatchTableSim#(25, 54, 26);
  function ActionValue#(Bit#(26)) matchtable_read(Bit#(25) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_ipv4_dest_vtep(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(25) id, Bit#(54) key, Bit#(26) data);
    action
      matchtable_write_ipv4_dest_vtep(key, data);
    endaction
  endfunction

endinstance
interface Ipv4DestVtep;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIpv4DestVtep  (Ipv4DestVtep);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(25, 1024, SizeOf#(Ipv4DestVtepReqT), SizeOf#(Ipv4DestVtepRspT)) matchTable <- mkMatchTable("ipv4_dest_vtep.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv4$dstAddr = fromMaybe(?, meta.ipv4$dstAddr);
    let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
    Ipv4DestVtepReqT req = Ipv4DestVtepReqT {l3_metadata$vrf: l3_metadata$vrf,ipv4$dstAddr: ipv4$dstAddr,tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4DestVtepRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_TUNNEL_TERMINATION_FLAG: begin
          BBRequest req = tagged SetTunnelTerminationFlagReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_TUNNEL_VNI_AND_TERMINATION_FLAG: begin
          BBRequest req = tagged SetTunnelVniAndTerminationFlagReqT {pkt: pkt, runtime_tunnel_vni: resp.runtime_tunnel_vni};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4DestVtepNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetTunnelTerminationFlagRspT {pkt: .pkt, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate}: begin
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        MetadataResponse rsp = tagged Ipv4DestVtepSetTunnelTerminationFlagRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetTunnelVniAndTerminationFlagRspT {pkt: .pkt, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, tunnel_metadata$tunnel_vni: .tunnel_metadata$tunnel_vni}: begin
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.tunnel_metadata$tunnel_vni = tagged Valid tunnel_metadata$tunnel_vni;
        MetadataResponse rsp = tagged Ipv4DestVtepSetTunnelVniAndTerminationFlagRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== IPV4_FIB ======

typedef struct {
  Bit#(6) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
} Ipv4FibReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_FIB,
  ON_MISS,
  FIB_HIT_NEXTHOP,
  FIB_HIT_ECMP
} Ipv4FibActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4FibActionT _action;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} Ipv4FibRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_ipv4_fib(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_ipv4_fib(Bit#(54) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(15, 54, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(15) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_ipv4_fib(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(15) id, Bit#(54) key, Bit#(34) data);
    action
      matchtable_write_ipv4_fib(key, data);
    endaction
  endfunction

endinstance
interface Ipv4Fib;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIpv4Fib  (Ipv4Fib);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(15, 1024, SizeOf#(Ipv4FibReqT), SizeOf#(Ipv4FibRspT)) matchTable <- mkMatchTable("ipv4_fib.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    Ipv4FibReqT req = Ipv4FibReqT {l3_metadata$vrf: l3_metadata$vrf,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4FibRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        FIB_HIT_NEXTHOP: begin
          BBRequest req = tagged FibHitNexthopReqT {pkt: pkt, runtime_nexthop_index: resp.runtime_nexthop_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        FIB_HIT_ECMP: begin
          BBRequest req = tagged FibHitEcmpReqT {pkt: pkt, runtime_ecmp_index: resp.runtime_ecmp_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4FibOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FibHitNexthopRspT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        MetadataResponse rsp = tagged Ipv4FibFibHitNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FibHitEcmpRspT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        MetadataResponse rsp = tagged Ipv4FibFibHitEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== IPV4_FIB_LPM ======

typedef struct {
  Bit#(6) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
} Ipv4FibLpmReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_FIB_LPM,
  ON_MISS,
  FIB_HIT_NEXTHOP,
  FIB_HIT_ECMP
} Ipv4FibLpmActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4FibLpmActionT _action;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} Ipv4FibLpmRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_ipv4_fib_lpm(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_ipv4_fib_lpm(Bit#(54) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(16, 54, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(16) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_ipv4_fib_lpm(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(16) id, Bit#(54) key, Bit#(34) data);
    action
      matchtable_write_ipv4_fib_lpm(key, data);
    endaction
  endfunction

endinstance
interface Ipv4FibLpm;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIpv4FibLpm  (Ipv4FibLpm);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(16, 512, SizeOf#(Ipv4FibLpmReqT), SizeOf#(Ipv4FibLpmRspT)) matchTable <- mkMatchTable("ipv4_fib_lpm.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    Ipv4FibLpmReqT req = Ipv4FibLpmReqT {l3_metadata$vrf: l3_metadata$vrf,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4FibLpmRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        FIB_HIT_NEXTHOP: begin
          BBRequest req = tagged FibHitNexthopReqT {pkt: pkt, runtime_nexthop_index: resp.runtime_nexthop_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        FIB_HIT_ECMP: begin
          BBRequest req = tagged FibHitEcmpReqT {pkt: pkt, runtime_ecmp_index: resp.runtime_ecmp_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4FibLpmOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FibHitNexthopRspT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        MetadataResponse rsp = tagged Ipv4FibLpmFibHitNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FibHitEcmpRspT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        MetadataResponse rsp = tagged Ipv4FibLpmFibHitEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== IPV4_MULTICAST_BRIDGE ======

typedef struct {
  Bit#(1) padding;
  Bit#(16) ingress_metadata$bd;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
} Ipv4MulticastBridgeReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_MULTICAST_BRIDGE,
  ON_MISS,
  MULTICAST_BRIDGE_S_G_HIT
} Ipv4MulticastBridgeActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4MulticastBridgeActionT _action;
  Bit#(16) runtime_mc_index;
} Ipv4MulticastBridgeRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv4_multicast_bridge(Bit#(81) msgtype);
import "BDPI" function Action matchtable_write_ipv4_multicast_bridge(Bit#(81) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(48, 81, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(48) id, Bit#(81) key);
    actionvalue
      let v <- matchtable_read_ipv4_multicast_bridge(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(48) id, Bit#(81) key, Bit#(18) data);
    action
      matchtable_write_ipv4_multicast_bridge(key, data);
    endaction
  endfunction

endinstance
interface Ipv4MulticastBridge;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv4MulticastBridge  (Ipv4MulticastBridge);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(48, 1024, SizeOf#(Ipv4MulticastBridgeReqT), SizeOf#(Ipv4MulticastBridgeRspT)) matchTable <- mkMatchTable("ipv4_multicast_bridge.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    Ipv4MulticastBridgeReqT req = Ipv4MulticastBridgeReqT {ingress_metadata$bd: ingress_metadata$bd,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4MulticastBridgeRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_BRIDGE_S_G_HIT: begin
          BBRequest req = tagged MulticastBridgeSGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4MulticastBridgeOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastBridgeSGHitRspT {pkt: .pkt, multicast_metadata$mcast_bridge_hit: .multicast_metadata$mcast_bridge_hit, multicast_metadata$multicast_bridge_mc_index: .multicast_metadata$multicast_bridge_mc_index}: begin
        meta.multicast_metadata$mcast_bridge_hit = tagged Valid multicast_metadata$mcast_bridge_hit;
        meta.multicast_metadata$multicast_bridge_mc_index = tagged Valid multicast_metadata$multicast_bridge_mc_index;
        MetadataResponse rsp = tagged Ipv4MulticastBridgeMulticastBridgeSGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV4_MULTICAST_BRIDGE_STAR_G ======

typedef struct {
  Bit#(6) padding;
  Bit#(16) ingress_metadata$bd;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
} Ipv4MulticastBridgeStarGReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_MULTICAST_BRIDGE_STAR_G,
  NOP,
  MULTICAST_BRIDGE_STAR_G_HIT
} Ipv4MulticastBridgeStarGActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4MulticastBridgeStarGActionT _action;
  Bit#(16) runtime_mc_index;
} Ipv4MulticastBridgeStarGRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv4_multicast_bridge_star_g(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_ipv4_multicast_bridge_star_g(Bit#(54) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(47, 54, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(47) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_ipv4_multicast_bridge_star_g(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(47) id, Bit#(54) key, Bit#(18) data);
    action
      matchtable_write_ipv4_multicast_bridge_star_g(key, data);
    endaction
  endfunction

endinstance
interface Ipv4MulticastBridgeStarG;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv4MulticastBridgeStarG  (Ipv4MulticastBridgeStarG);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(47, 1024, SizeOf#(Ipv4MulticastBridgeStarGReqT), SizeOf#(Ipv4MulticastBridgeStarGRspT)) matchTable <- mkMatchTable("ipv4_multicast_bridge_star_g.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    Ipv4MulticastBridgeStarGReqT req = Ipv4MulticastBridgeStarGReqT {ingress_metadata$bd: ingress_metadata$bd,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4MulticastBridgeStarGRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_BRIDGE_STAR_G_HIT: begin
          BBRequest req = tagged MulticastBridgeStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4MulticastBridgeStarGNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastBridgeStarGHitRspT {pkt: .pkt, multicast_metadata$mcast_bridge_hit: .multicast_metadata$mcast_bridge_hit, multicast_metadata$multicast_bridge_mc_index: .multicast_metadata$multicast_bridge_mc_index}: begin
        meta.multicast_metadata$mcast_bridge_hit = tagged Valid multicast_metadata$mcast_bridge_hit;
        meta.multicast_metadata$multicast_bridge_mc_index = tagged Valid multicast_metadata$multicast_bridge_mc_index;
        MetadataResponse rsp = tagged Ipv4MulticastBridgeStarGMulticastBridgeStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV4_MULTICAST_ROUTE ======

typedef struct {
  Bit#(1) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
} Ipv4MulticastRouteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_MULTICAST_ROUTE,
  ON_MISS,
  MULTICAST_ROUTE_S_G_HIT
} Ipv4MulticastRouteActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4MulticastRouteActionT _action;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_mcast_rpf_group;
} Ipv4MulticastRouteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_ipv4_multicast_route(Bit#(81) msgtype);
import "BDPI" function Action matchtable_write_ipv4_multicast_route(Bit#(81) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(50, 81, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(50) id, Bit#(81) key);
    actionvalue
      let v <- matchtable_read_ipv4_multicast_route(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(50) id, Bit#(81) key, Bit#(34) data);
    action
      matchtable_write_ipv4_multicast_route(key, data);
    endaction
  endfunction

endinstance
interface Ipv4MulticastRoute;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv4MulticastRoute  (Ipv4MulticastRoute);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(50, 1024, SizeOf#(Ipv4MulticastRouteReqT), SizeOf#(Ipv4MulticastRouteRspT)) matchTable <- mkMatchTable("ipv4_multicast_route.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    Ipv4MulticastRouteReqT req = Ipv4MulticastRouteReqT {l3_metadata$vrf: l3_metadata$vrf,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4MulticastRouteRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_ROUTE_S_G_HIT: begin
          BBRequest req = tagged MulticastRouteSGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4MulticastRouteOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastRouteSGHitRspT {pkt: .pkt, multicast_metadata$mcast_route_hit: .multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: .multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: .multicast_metadata$mcast_mode}: begin
        meta.multicast_metadata$mcast_route_hit = tagged Valid multicast_metadata$mcast_route_hit;
        meta.multicast_metadata$multicast_route_mc_index = tagged Valid multicast_metadata$multicast_route_mc_index;
        meta.multicast_metadata$mcast_mode = tagged Valid multicast_metadata$mcast_mode;
        MetadataResponse rsp = tagged Ipv4MulticastRouteMulticastRouteSGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV4_MULTICAST_ROUTE_STAR_G ======

typedef struct {
  Bit#(6) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
} Ipv4MulticastRouteStarGReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_MULTICAST_ROUTE_STAR_G,
  MULTICAST_ROUTE_STAR_G_MISS,
  MULTICAST_ROUTE_SM_STAR_G_HIT,
  MULTICAST_ROUTE_BIDIR_STAR_G_HIT
} Ipv4MulticastRouteStarGActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4MulticastRouteStarGActionT _action;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_mcast_rpf_group;
} Ipv4MulticastRouteStarGRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_ipv4_multicast_route_star_g(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_ipv4_multicast_route_star_g(Bit#(54) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(49, 54, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(49) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_ipv4_multicast_route_star_g(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(49) id, Bit#(54) key, Bit#(34) data);
    action
      matchtable_write_ipv4_multicast_route_star_g(key, data);
    endaction
  endfunction

endinstance
interface Ipv4MulticastRouteStarG;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIpv4MulticastRouteStarG  (Ipv4MulticastRouteStarG);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(49, 1024, SizeOf#(Ipv4MulticastRouteStarGReqT), SizeOf#(Ipv4MulticastRouteStarGRspT)) matchTable <- mkMatchTable("ipv4_multicast_route_star_g.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    Ipv4MulticastRouteStarGReqT req = Ipv4MulticastRouteStarGReqT {l3_metadata$vrf: l3_metadata$vrf,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4MulticastRouteStarGRspT resp = unpack(data);
      case (resp._action) matches
        MULTICAST_ROUTE_STAR_G_MISS: begin
          BBRequest req = tagged MulticastRouteStarGMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_ROUTE_SM_STAR_G_HIT: begin
          BBRequest req = tagged MulticastRouteSmStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_ROUTE_BIDIR_STAR_G_HIT: begin
          BBRequest req = tagged MulticastRouteBidirStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged MulticastRouteStarGMissRspT {pkt: .pkt, l3_metadata$l3_copy: .l3_metadata$l3_copy}: begin
        meta.l3_metadata$l3_copy = tagged Valid l3_metadata$l3_copy;
        MetadataResponse rsp = tagged Ipv4MulticastRouteStarGMulticastRouteStarGMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastRouteSmStarGHitRspT {pkt: .pkt, multicast_metadata$mcast_route_hit: .multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: .multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: .multicast_metadata$mcast_mode}: begin
        meta.multicast_metadata$mcast_route_hit = tagged Valid multicast_metadata$mcast_route_hit;
        meta.multicast_metadata$multicast_route_mc_index = tagged Valid multicast_metadata$multicast_route_mc_index;
        meta.multicast_metadata$mcast_mode = tagged Valid multicast_metadata$mcast_mode;
        MetadataResponse rsp = tagged Ipv4MulticastRouteStarGMulticastRouteSmStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastRouteBidirStarGHitRspT {pkt: .pkt, multicast_metadata$mcast_route_hit: .multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: .multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: .multicast_metadata$mcast_mode}: begin
        meta.multicast_metadata$mcast_route_hit = tagged Valid multicast_metadata$mcast_route_hit;
        meta.multicast_metadata$multicast_route_mc_index = tagged Valid multicast_metadata$multicast_route_mc_index;
        meta.multicast_metadata$mcast_mode = tagged Valid multicast_metadata$mcast_mode;
        MetadataResponse rsp = tagged Ipv4MulticastRouteStarGMulticastRouteBidirStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== IPV4_RACL ======

typedef struct {
  Bit#(6) padding;
  Bit#(16) acl_metadata$bd_label;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
  Bit#(8) l3_metadata$lkp_ip_proto;
  Bit#(16) l3_metadata$lkp_l4_sport;
  Bit#(16) l3_metadata$lkp_l4_dport;
} Ipv4RaclReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_RACL,
  NOP,
  RACL_DENY,
  RACL_PERMIT,
  RACL_REDIRECT_NEXTHOP,
  RACL_REDIRECT_ECMP
} Ipv4RaclActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4RaclActionT _action;
  Bit#(14) runtime_acl_stats_index;
  Bit#(1) runtime_acl_copy;
  Bit#(16) runtime_acl_copy_reason;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} Ipv4RaclRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(66)) matchtable_read_ipv4_racl(Bit#(126) msgtype);
import "BDPI" function Action matchtable_write_ipv4_racl(Bit#(126) msgtype, Bit#(66) data);
`endif
instance MatchTableSim#(38, 126, 66);
  function ActionValue#(Bit#(66)) matchtable_read(Bit#(38) id, Bit#(126) key);
    actionvalue
      let v <- matchtable_read_ipv4_racl(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(38) id, Bit#(126) key, Bit#(66) data);
    action
      matchtable_write_ipv4_racl(key, data);
    endaction
  endfunction

endinstance
interface Ipv4Racl;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
endinterface
(* synthesize *)
module mkIpv4Racl  (Ipv4Racl);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(5, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(5, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(38, 512, SizeOf#(Ipv4RaclReqT), SizeOf#(Ipv4RaclRspT)) matchTable <- mkMatchTable("ipv4_racl.dat");
  Vector#(5, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(5) readyChannel = -1;
  for (Integer i=4; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let acl_metadata$bd_label = fromMaybe(?, meta.acl_metadata$bd_label);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    let l3_metadata$lkp_ip_proto = fromMaybe(?, meta.l3_metadata$lkp_ip_proto);
    let l3_metadata$lkp_l4_sport = fromMaybe(?, meta.l3_metadata$lkp_l4_sport);
    let l3_metadata$lkp_l4_dport = fromMaybe(?, meta.l3_metadata$lkp_l4_dport);
    Ipv4RaclReqT req = Ipv4RaclReqT {acl_metadata$bd_label: acl_metadata$bd_label,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da,l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto,l3_metadata$lkp_l4_sport: l3_metadata$lkp_l4_sport,l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4RaclRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        RACL_DENY: begin
          BBRequest req = tagged RaclDenyReqT {pkt: pkt, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        RACL_PERMIT: begin
          BBRequest req = tagged RaclPermitReqT {pkt: pkt, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        RACL_REDIRECT_NEXTHOP: begin
          BBRequest req = tagged RaclRedirectNexthopReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_nexthop_index: resp.runtime_nexthop_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        RACL_REDIRECT_ECMP: begin
          BBRequest req = tagged RaclRedirectEcmpReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_ecmp_index: resp.runtime_ecmp_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4RaclNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RaclDenyRspT {pkt: .pkt, acl_metadata$racl_deny: .acl_metadata$racl_deny, acl_metadata$acl_copy: .acl_metadata$acl_copy, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index}: begin
        meta.acl_metadata$racl_deny = tagged Valid acl_metadata$racl_deny;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        MetadataResponse rsp = tagged Ipv4RaclRaclDenyRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RaclPermitRspT {pkt: .pkt, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$acl_copy: .acl_metadata$acl_copy, fabric_metadata$reason_code: .fabric_metadata$reason_code}: begin
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        MetadataResponse rsp = tagged Ipv4RaclRaclPermitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RaclRedirectNexthopRspT {pkt: .pkt, acl_metadata$racl_nexthop: .acl_metadata$racl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$racl_redirect: .acl_metadata$racl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$racl_nexthop_type: .acl_metadata$racl_nexthop_type}: begin
        meta.acl_metadata$racl_nexthop = tagged Valid acl_metadata$racl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$racl_redirect = tagged Valid acl_metadata$racl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$racl_nexthop_type = tagged Valid acl_metadata$racl_nexthop_type;
        MetadataResponse rsp = tagged Ipv4RaclRaclRedirectNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RaclRedirectEcmpRspT {pkt: .pkt, acl_metadata$racl_nexthop: .acl_metadata$racl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$racl_redirect: .acl_metadata$racl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$racl_nexthop_type: .acl_metadata$racl_nexthop_type}: begin
        meta.acl_metadata$racl_nexthop = tagged Valid acl_metadata$racl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$racl_redirect = tagged Valid acl_metadata$racl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$racl_nexthop_type = tagged Valid acl_metadata$racl_nexthop_type;
        MetadataResponse rsp = tagged Ipv4RaclRaclRedirectEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
endmodule

// ====== IPV4_SRC_VTEP ======

typedef struct {
  Bit#(1) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(32) ipv4$srcAddr;
  Bit#(5) tunnel_metadata$ingress_tunnel_type;
} Ipv4SrcVtepReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_SRC_VTEP,
  ON_MISS,
  SRC_VTEP_HIT
} Ipv4SrcVtepActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4SrcVtepActionT _action;
  Bit#(16) runtime_ifindex;
} Ipv4SrcVtepRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv4_src_vtep(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_ipv4_src_vtep(Bit#(54) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(26, 54, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(26) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_ipv4_src_vtep(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(26) id, Bit#(54) key, Bit#(18) data);
    action
      matchtable_write_ipv4_src_vtep(key, data);
    endaction
  endfunction

endinstance
interface Ipv4SrcVtep;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv4SrcVtep  (Ipv4SrcVtep);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(26, 1024, SizeOf#(Ipv4SrcVtepReqT), SizeOf#(Ipv4SrcVtepRspT)) matchTable <- mkMatchTable("ipv4_src_vtep.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv4$srcAddr = fromMaybe(?, meta.ipv4$srcAddr);
    let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
    Ipv4SrcVtepReqT req = Ipv4SrcVtepReqT {l3_metadata$vrf: l3_metadata$vrf,ipv4$srcAddr: ipv4$srcAddr,tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4SrcVtepRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SRC_VTEP_HIT: begin
          BBRequest req = tagged SrcVtepHitReqT {pkt: pkt, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4SrcVtepOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SrcVtepHitRspT {pkt: .pkt, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        meta.ingress_metadata$ifindex = tagged Valid ingress_metadata$ifindex;
        MetadataResponse rsp = tagged Ipv4SrcVtepSrcVtepHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV4_URPF ======

typedef struct {
  Bit#(6) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
} Ipv4UrpfReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_URPF,
  ON_MISS,
  IPV4_URPF_HIT
} Ipv4UrpfActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4UrpfActionT _action;
  Bit#(16) runtime_urpf_bd_group;
} Ipv4UrpfRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv4_urpf(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_ipv4_urpf(Bit#(54) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(18, 54, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(18) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_ipv4_urpf(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(18) id, Bit#(54) key, Bit#(18) data);
    action
      matchtable_write_ipv4_urpf(key, data);
    endaction
  endfunction

endinstance
interface Ipv4Urpf;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv4Urpf  (Ipv4Urpf);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(18, 1024, SizeOf#(Ipv4UrpfReqT), SizeOf#(Ipv4UrpfRspT)) matchTable <- mkMatchTable("ipv4_urpf.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    Ipv4UrpfReqT req = Ipv4UrpfReqT {l3_metadata$vrf: l3_metadata$vrf,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4UrpfRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_URPF_HIT: begin
          BBRequest req = tagged Ipv4UrpfHitReqT {pkt: pkt, ipv4_metadata$ipv4_urpf_mode: ipv4_metadata$ipv4_urpf_mode, runtime_urpf_bd_group: resp.runtime_urpf_bd_group};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv4UrpfOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4UrpfHitRspT {pkt: .pkt, l3_metadata$urpf_bd_group: .l3_metadata$urpf_bd_group, l3_metadata$urpf_hit: .l3_metadata$urpf_hit, l3_metadata$urpf_mode: .l3_metadata$urpf_mode}: begin
        meta.l3_metadata$urpf_bd_group = tagged Valid l3_metadata$urpf_bd_group;
        meta.l3_metadata$urpf_hit = tagged Valid l3_metadata$urpf_hit;
        meta.l3_metadata$urpf_mode = tagged Valid l3_metadata$urpf_mode;
        MetadataResponse rsp = tagged Ipv4UrpfIpv4UrpfHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV4_URPF_LPM ======

typedef struct {
  Bit#(6) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
} Ipv4UrpfLpmReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV4_URPF_LPM,
  IPV4_URPF_HIT,
  URPF_MISS
} Ipv4UrpfLpmActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv4UrpfLpmActionT _action;
  Bit#(16) runtime_urpf_bd_group;
} Ipv4UrpfLpmRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv4_urpf_lpm(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_ipv4_urpf_lpm(Bit#(54) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(17, 54, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(17) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_ipv4_urpf_lpm(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(17) id, Bit#(54) key, Bit#(18) data);
    action
      matchtable_write_ipv4_urpf_lpm(key, data);
    endaction
  endfunction

endinstance
interface Ipv4UrpfLpm;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv4UrpfLpm  (Ipv4UrpfLpm);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(17, 512, SizeOf#(Ipv4UrpfLpmReqT), SizeOf#(Ipv4UrpfLpmRspT)) matchTable <- mkMatchTable("ipv4_urpf_lpm.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    Ipv4UrpfLpmReqT req = Ipv4UrpfLpmReqT {l3_metadata$vrf: l3_metadata$vrf,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv4UrpfLpmRspT resp = unpack(data);
      case (resp._action) matches
        IPV4_URPF_HIT: begin
          BBRequest req = tagged Ipv4UrpfHitReqT {pkt: pkt, ipv4_metadata$ipv4_urpf_mode: ipv4_metadata$ipv4_urpf_mode, runtime_urpf_bd_group: resp.runtime_urpf_bd_group};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        URPF_MISS: begin
          BBRequest req = tagged UrpfMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged Ipv4UrpfHitRspT {pkt: .pkt, l3_metadata$urpf_bd_group: .l3_metadata$urpf_bd_group, l3_metadata$urpf_hit: .l3_metadata$urpf_hit, l3_metadata$urpf_mode: .l3_metadata$urpf_mode}: begin
        meta.l3_metadata$urpf_bd_group = tagged Valid l3_metadata$urpf_bd_group;
        meta.l3_metadata$urpf_hit = tagged Valid l3_metadata$urpf_hit;
        meta.l3_metadata$urpf_mode = tagged Valid l3_metadata$urpf_mode;
        MetadataResponse rsp = tagged Ipv4UrpfLpmIpv4UrpfHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged UrpfMissRspT {pkt: .pkt, l3_metadata$urpf_check_fail: .l3_metadata$urpf_check_fail}: begin
        meta.l3_metadata$urpf_check_fail = tagged Valid l3_metadata$urpf_check_fail;
        MetadataResponse rsp = tagged Ipv4UrpfLpmUrpfMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV6_ACL ======

typedef struct {
  Bit#(7) padding;
  Bit#(16) acl_metadata$if_label;
  Bit#(16) acl_metadata$bd_label;
  Bit#(128) ipv6_metadata$lkp_ipv6_sa;
  Bit#(128) ipv6_metadata$lkp_ipv6_da;
  Bit#(8) l3_metadata$lkp_ip_proto;
  Bit#(16) l3_metadata$lkp_l4_sport;
  Bit#(16) l3_metadata$lkp_l4_dport;
  Bit#(8) tcp$flags;
  Bit#(8) l3_metadata$lkp_ip_ttl;
} Ipv6AclReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_ACL,
  NOP,
  ACL_DENY,
  ACL_PERMIT,
  ACL_MIRROR,
  ACL_REDIRECT_NEXTHOP,
  ACL_REDIRECT_ECMP
} Ipv6AclActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6AclActionT _action;
  Bit#(14) runtime_acl_stats_index;
  Bit#(16) runtime_acl_meter_index;
  Bit#(1) runtime_acl_copy;
  Bit#(16) runtime_acl_copy_reason;
  Bit#(32) runtime_session_id;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} Ipv6AclRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(114)) matchtable_read_ipv6_acl(Bit#(351) msgtype);
import "BDPI" function Action matchtable_write_ipv6_acl(Bit#(351) msgtype, Bit#(114) data);
`endif
instance MatchTableSim#(36, 351, 114);
  function ActionValue#(Bit#(114)) matchtable_read(Bit#(36) id, Bit#(351) key);
    actionvalue
      let v <- matchtable_read_ipv6_acl(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(36) id, Bit#(351) key, Bit#(114) data);
    action
      matchtable_write_ipv6_acl(key, data);
    endaction
  endfunction

endinstance
interface Ipv6Acl;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
endinterface
(* synthesize *)
module mkIpv6Acl  (Ipv6Acl);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(6, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(6, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(36, 512, SizeOf#(Ipv6AclReqT), SizeOf#(Ipv6AclRspT)) matchTable <- mkMatchTable("ipv6_acl.dat");
  Vector#(6, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(6) readyChannel = -1;
  for (Integer i=5; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let acl_metadata$if_label = fromMaybe(?, meta.acl_metadata$if_label);
    let acl_metadata$bd_label = fromMaybe(?, meta.acl_metadata$bd_label);
    let ipv6_metadata$lkp_ipv6_sa = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_sa);
    let ipv6_metadata$lkp_ipv6_da = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_da);
    let l3_metadata$lkp_ip_proto = fromMaybe(?, meta.l3_metadata$lkp_ip_proto);
    let l3_metadata$lkp_l4_sport = fromMaybe(?, meta.l3_metadata$lkp_l4_sport);
    let l3_metadata$lkp_l4_dport = fromMaybe(?, meta.l3_metadata$lkp_l4_dport);
    let tcp$flags = fromMaybe(?, meta.tcp$flags);
    let l3_metadata$lkp_ip_ttl = fromMaybe(?, meta.l3_metadata$lkp_ip_ttl);
    Ipv6AclReqT req = Ipv6AclReqT {acl_metadata$if_label: acl_metadata$if_label,acl_metadata$bd_label: acl_metadata$bd_label,ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa,ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da,l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto,l3_metadata$lkp_l4_sport: l3_metadata$lkp_l4_sport,l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport,tcp$flags: tcp$flags,l3_metadata$lkp_ip_ttl: l3_metadata$lkp_ip_ttl};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6AclRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        ACL_DENY: begin
          BBRequest req = tagged AclDenyReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        ACL_PERMIT: begin
          BBRequest req = tagged AclPermitReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        ACL_MIRROR: begin
          BBRequest req = tagged AclMirrorReqT {pkt: pkt, intrinsic_metadata$ingress_global_tstamp: intrinsic_metadata$ingress_global_tstamp, runtime_session_id: resp.runtime_session_id, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        ACL_REDIRECT_NEXTHOP: begin
          BBRequest req = tagged AclRedirectNexthopReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_copy: resp.runtime_acl_copy, runtime_nexthop_index: resp.runtime_nexthop_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        ACL_REDIRECT_ECMP: begin
          BBRequest req = tagged AclRedirectEcmpReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_copy: resp.runtime_acl_copy, runtime_ecmp_index: resp.runtime_ecmp_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6AclNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclDenyRspT {pkt: .pkt, acl_metadata$acl_deny: .acl_metadata$acl_deny, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_copy: .acl_metadata$acl_copy}: begin
        meta.acl_metadata$acl_deny = tagged Valid acl_metadata$acl_deny;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        MetadataResponse rsp = tagged Ipv6AclAclDenyRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclPermitRspT {pkt: .pkt, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_copy: .acl_metadata$acl_copy}: begin
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        MetadataResponse rsp = tagged Ipv6AclAclPermitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclMirrorRspT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id}: begin
        meta.i2e_metadata$ingress_tstamp = tagged Valid i2e_metadata$ingress_tstamp;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.i2e_metadata$mirror_session_id = tagged Valid i2e_metadata$mirror_session_id;
        MetadataResponse rsp = tagged Ipv6AclAclMirrorRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclRedirectNexthopRspT {pkt: .pkt, meter_metadata$meter_index: .meter_metadata$meter_index, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$acl_redirect: .acl_metadata$acl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_nexthop: .acl_metadata$acl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_nexthop_type: .acl_metadata$acl_nexthop_type}: begin
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$acl_redirect = tagged Valid acl_metadata$acl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_nexthop = tagged Valid acl_metadata$acl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_nexthop_type = tagged Valid acl_metadata$acl_nexthop_type;
        MetadataResponse rsp = tagged Ipv6AclAclRedirectNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclRedirectEcmpRspT {pkt: .pkt, meter_metadata$meter_index: .meter_metadata$meter_index, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$acl_redirect: .acl_metadata$acl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_nexthop: .acl_metadata$acl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_nexthop_type: .acl_metadata$acl_nexthop_type}: begin
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$acl_redirect = tagged Valid acl_metadata$acl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_nexthop = tagged Valid acl_metadata$acl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_nexthop_type = tagged Valid acl_metadata$acl_nexthop_type;
        MetadataResponse rsp = tagged Ipv6AclAclRedirectEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
endmodule

// ====== IPV6_DEST_VTEP ======

typedef struct {
  Bit#(4) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(128) ipv6$dstAddr;
  Bit#(5) tunnel_metadata$ingress_tunnel_type;
} Ipv6DestVtepReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_DEST_VTEP,
  NOP,
  SET_TUNNEL_TERMINATION_FLAG,
  SET_TUNNEL_VNI_AND_TERMINATION_FLAG
} Ipv6DestVtepActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6DestVtepActionT _action;
  Bit#(24) runtime_tunnel_vni;
} Ipv6DestVtepRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(26)) matchtable_read_ipv6_dest_vtep(Bit#(153) msgtype);
import "BDPI" function Action matchtable_write_ipv6_dest_vtep(Bit#(153) msgtype, Bit#(26) data);
`endif
instance MatchTableSim#(27, 153, 26);
  function ActionValue#(Bit#(26)) matchtable_read(Bit#(27) id, Bit#(153) key);
    actionvalue
      let v <- matchtable_read_ipv6_dest_vtep(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(27) id, Bit#(153) key, Bit#(26) data);
    action
      matchtable_write_ipv6_dest_vtep(key, data);
    endaction
  endfunction

endinstance
interface Ipv6DestVtep;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIpv6DestVtep  (Ipv6DestVtep);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(27, 1024, SizeOf#(Ipv6DestVtepReqT), SizeOf#(Ipv6DestVtepRspT)) matchTable <- mkMatchTable("ipv6_dest_vtep.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv6$dstAddr = fromMaybe(?, meta.ipv6$dstAddr);
    let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
    Ipv6DestVtepReqT req = Ipv6DestVtepReqT {l3_metadata$vrf: l3_metadata$vrf,ipv6$dstAddr: ipv6$dstAddr,tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6DestVtepRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_TUNNEL_TERMINATION_FLAG: begin
          BBRequest req = tagged SetTunnelTerminationFlagReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_TUNNEL_VNI_AND_TERMINATION_FLAG: begin
          BBRequest req = tagged SetTunnelVniAndTerminationFlagReqT {pkt: pkt, runtime_tunnel_vni: resp.runtime_tunnel_vni};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6DestVtepNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetTunnelTerminationFlagRspT {pkt: .pkt, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate}: begin
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        MetadataResponse rsp = tagged Ipv6DestVtepSetTunnelTerminationFlagRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetTunnelVniAndTerminationFlagRspT {pkt: .pkt, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, tunnel_metadata$tunnel_vni: .tunnel_metadata$tunnel_vni}: begin
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.tunnel_metadata$tunnel_vni = tagged Valid tunnel_metadata$tunnel_vni;
        MetadataResponse rsp = tagged Ipv6DestVtepSetTunnelVniAndTerminationFlagRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== IPV6_FIB ======

typedef struct {
  Bit#(16) l3_metadata$vrf;
  Bit#(128) ipv6_metadata$lkp_ipv6_da;
} Ipv6FibReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_FIB,
  ON_MISS,
  FIB_HIT_NEXTHOP,
  FIB_HIT_ECMP
} Ipv6FibActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6FibActionT _action;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} Ipv6FibRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_ipv6_fib(Bit#(144) msgtype);
import "BDPI" function Action matchtable_write_ipv6_fib(Bit#(144) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(21, 144, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(21) id, Bit#(144) key);
    actionvalue
      let v <- matchtable_read_ipv6_fib(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(21) id, Bit#(144) key, Bit#(34) data);
    action
      matchtable_write_ipv6_fib(key, data);
    endaction
  endfunction

endinstance
interface Ipv6Fib;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIpv6Fib  (Ipv6Fib);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(21, 1024, SizeOf#(Ipv6FibReqT), SizeOf#(Ipv6FibRspT)) matchTable <- mkMatchTable("ipv6_fib.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv6_metadata$lkp_ipv6_da = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_da);
    Ipv6FibReqT req = Ipv6FibReqT {l3_metadata$vrf: l3_metadata$vrf,ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6FibRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        FIB_HIT_NEXTHOP: begin
          BBRequest req = tagged FibHitNexthopReqT {pkt: pkt, runtime_nexthop_index: resp.runtime_nexthop_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        FIB_HIT_ECMP: begin
          BBRequest req = tagged FibHitEcmpReqT {pkt: pkt, runtime_ecmp_index: resp.runtime_ecmp_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6FibOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FibHitNexthopRspT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        MetadataResponse rsp = tagged Ipv6FibFibHitNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FibHitEcmpRspT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        MetadataResponse rsp = tagged Ipv6FibFibHitEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== IPV6_FIB_LPM ======

typedef struct {
  Bit#(16) l3_metadata$vrf;
  Bit#(128) ipv6_metadata$lkp_ipv6_da;
} Ipv6FibLpmReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_FIB_LPM,
  ON_MISS,
  FIB_HIT_NEXTHOP,
  FIB_HIT_ECMP
} Ipv6FibLpmActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6FibLpmActionT _action;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} Ipv6FibLpmRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_ipv6_fib_lpm(Bit#(144) msgtype);
import "BDPI" function Action matchtable_write_ipv6_fib_lpm(Bit#(144) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(20, 144, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(20) id, Bit#(144) key);
    actionvalue
      let v <- matchtable_read_ipv6_fib_lpm(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(20) id, Bit#(144) key, Bit#(34) data);
    action
      matchtable_write_ipv6_fib_lpm(key, data);
    endaction
  endfunction

endinstance
interface Ipv6FibLpm;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIpv6FibLpm  (Ipv6FibLpm);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(20, 512, SizeOf#(Ipv6FibLpmReqT), SizeOf#(Ipv6FibLpmRspT)) matchTable <- mkMatchTable("ipv6_fib_lpm.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv6_metadata$lkp_ipv6_da = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_da);
    Ipv6FibLpmReqT req = Ipv6FibLpmReqT {l3_metadata$vrf: l3_metadata$vrf,ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6FibLpmRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        FIB_HIT_NEXTHOP: begin
          BBRequest req = tagged FibHitNexthopReqT {pkt: pkt, runtime_nexthop_index: resp.runtime_nexthop_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        FIB_HIT_ECMP: begin
          BBRequest req = tagged FibHitEcmpReqT {pkt: pkt, runtime_ecmp_index: resp.runtime_ecmp_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6FibLpmOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FibHitNexthopRspT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        MetadataResponse rsp = tagged Ipv6FibLpmFibHitNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FibHitEcmpRspT {pkt: .pkt, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type}: begin
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        MetadataResponse rsp = tagged Ipv6FibLpmFibHitEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== IPV6_MULTICAST_BRIDGE ======

typedef struct {
  Bit#(7) padding;
  Bit#(16) ingress_metadata$bd;
  Bit#(128) ipv6_metadata$lkp_ipv6_sa;
  Bit#(128) ipv6_metadata$lkp_ipv6_da;
} Ipv6MulticastBridgeReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_MULTICAST_BRIDGE,
  ON_MISS,
  MULTICAST_BRIDGE_S_G_HIT
} Ipv6MulticastBridgeActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6MulticastBridgeActionT _action;
  Bit#(16) runtime_mc_index;
} Ipv6MulticastBridgeRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv6_multicast_bridge(Bit#(279) msgtype);
import "BDPI" function Action matchtable_write_ipv6_multicast_bridge(Bit#(279) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(52, 279, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(52) id, Bit#(279) key);
    actionvalue
      let v <- matchtable_read_ipv6_multicast_bridge(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(52) id, Bit#(279) key, Bit#(18) data);
    action
      matchtable_write_ipv6_multicast_bridge(key, data);
    endaction
  endfunction

endinstance
interface Ipv6MulticastBridge;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv6MulticastBridge  (Ipv6MulticastBridge);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(52, 1024, SizeOf#(Ipv6MulticastBridgeReqT), SizeOf#(Ipv6MulticastBridgeRspT)) matchTable <- mkMatchTable("ipv6_multicast_bridge.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    let ipv6_metadata$lkp_ipv6_sa = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_sa);
    let ipv6_metadata$lkp_ipv6_da = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_da);
    Ipv6MulticastBridgeReqT req = Ipv6MulticastBridgeReqT {ingress_metadata$bd: ingress_metadata$bd,ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa,ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6MulticastBridgeRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_BRIDGE_S_G_HIT: begin
          BBRequest req = tagged MulticastBridgeSGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6MulticastBridgeOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastBridgeSGHitRspT {pkt: .pkt, multicast_metadata$mcast_bridge_hit: .multicast_metadata$mcast_bridge_hit, multicast_metadata$multicast_bridge_mc_index: .multicast_metadata$multicast_bridge_mc_index}: begin
        meta.multicast_metadata$mcast_bridge_hit = tagged Valid multicast_metadata$mcast_bridge_hit;
        meta.multicast_metadata$multicast_bridge_mc_index = tagged Valid multicast_metadata$multicast_bridge_mc_index;
        MetadataResponse rsp = tagged Ipv6MulticastBridgeMulticastBridgeSGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV6_MULTICAST_BRIDGE_STAR_G ======

typedef struct {
  Bit#(16) ingress_metadata$bd;
  Bit#(128) ipv6_metadata$lkp_ipv6_da;
} Ipv6MulticastBridgeStarGReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_MULTICAST_BRIDGE_STAR_G,
  NOP,
  MULTICAST_BRIDGE_STAR_G_HIT
} Ipv6MulticastBridgeStarGActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6MulticastBridgeStarGActionT _action;
  Bit#(16) runtime_mc_index;
} Ipv6MulticastBridgeStarGRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv6_multicast_bridge_star_g(Bit#(144) msgtype);
import "BDPI" function Action matchtable_write_ipv6_multicast_bridge_star_g(Bit#(144) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(51, 144, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(51) id, Bit#(144) key);
    actionvalue
      let v <- matchtable_read_ipv6_multicast_bridge_star_g(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(51) id, Bit#(144) key, Bit#(18) data);
    action
      matchtable_write_ipv6_multicast_bridge_star_g(key, data);
    endaction
  endfunction

endinstance
interface Ipv6MulticastBridgeStarG;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv6MulticastBridgeStarG  (Ipv6MulticastBridgeStarG);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(51, 1024, SizeOf#(Ipv6MulticastBridgeStarGReqT), SizeOf#(Ipv6MulticastBridgeStarGRspT)) matchTable <- mkMatchTable("ipv6_multicast_bridge_star_g.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    let ipv6_metadata$lkp_ipv6_da = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_da);
    Ipv6MulticastBridgeStarGReqT req = Ipv6MulticastBridgeStarGReqT {ingress_metadata$bd: ingress_metadata$bd,ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6MulticastBridgeStarGRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_BRIDGE_STAR_G_HIT: begin
          BBRequest req = tagged MulticastBridgeStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6MulticastBridgeStarGNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastBridgeStarGHitRspT {pkt: .pkt, multicast_metadata$mcast_bridge_hit: .multicast_metadata$mcast_bridge_hit, multicast_metadata$multicast_bridge_mc_index: .multicast_metadata$multicast_bridge_mc_index}: begin
        meta.multicast_metadata$mcast_bridge_hit = tagged Valid multicast_metadata$mcast_bridge_hit;
        meta.multicast_metadata$multicast_bridge_mc_index = tagged Valid multicast_metadata$multicast_bridge_mc_index;
        MetadataResponse rsp = tagged Ipv6MulticastBridgeStarGMulticastBridgeStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV6_MULTICAST_ROUTE ======

typedef struct {
  Bit#(7) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(128) ipv6_metadata$lkp_ipv6_sa;
  Bit#(128) ipv6_metadata$lkp_ipv6_da;
} Ipv6MulticastRouteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_MULTICAST_ROUTE,
  ON_MISS,
  MULTICAST_ROUTE_S_G_HIT
} Ipv6MulticastRouteActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6MulticastRouteActionT _action;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_mcast_rpf_group;
} Ipv6MulticastRouteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_ipv6_multicast_route(Bit#(279) msgtype);
import "BDPI" function Action matchtable_write_ipv6_multicast_route(Bit#(279) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(54, 279, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(54) id, Bit#(279) key);
    actionvalue
      let v <- matchtable_read_ipv6_multicast_route(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(54) id, Bit#(279) key, Bit#(34) data);
    action
      matchtable_write_ipv6_multicast_route(key, data);
    endaction
  endfunction

endinstance
interface Ipv6MulticastRoute;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv6MulticastRoute  (Ipv6MulticastRoute);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(54, 1024, SizeOf#(Ipv6MulticastRouteReqT), SizeOf#(Ipv6MulticastRouteRspT)) matchTable <- mkMatchTable("ipv6_multicast_route.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv6_metadata$lkp_ipv6_sa = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_sa);
    let ipv6_metadata$lkp_ipv6_da = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_da);
    Ipv6MulticastRouteReqT req = Ipv6MulticastRouteReqT {l3_metadata$vrf: l3_metadata$vrf,ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa,ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6MulticastRouteRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_ROUTE_S_G_HIT: begin
          BBRequest req = tagged MulticastRouteSGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6MulticastRouteOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastRouteSGHitRspT {pkt: .pkt, multicast_metadata$mcast_route_hit: .multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: .multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: .multicast_metadata$mcast_mode}: begin
        meta.multicast_metadata$mcast_route_hit = tagged Valid multicast_metadata$mcast_route_hit;
        meta.multicast_metadata$multicast_route_mc_index = tagged Valid multicast_metadata$multicast_route_mc_index;
        meta.multicast_metadata$mcast_mode = tagged Valid multicast_metadata$mcast_mode;
        MetadataResponse rsp = tagged Ipv6MulticastRouteMulticastRouteSGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV6_MULTICAST_ROUTE_STAR_G ======

typedef struct {
  Bit#(16) l3_metadata$vrf;
  Bit#(128) ipv6_metadata$lkp_ipv6_da;
} Ipv6MulticastRouteStarGReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_MULTICAST_ROUTE_STAR_G,
  MULTICAST_ROUTE_STAR_G_MISS,
  MULTICAST_ROUTE_SM_STAR_G_HIT,
  MULTICAST_ROUTE_BIDIR_STAR_G_HIT
} Ipv6MulticastRouteStarGActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6MulticastRouteStarGActionT _action;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_mcast_rpf_group;
} Ipv6MulticastRouteStarGRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_ipv6_multicast_route_star_g(Bit#(144) msgtype);
import "BDPI" function Action matchtable_write_ipv6_multicast_route_star_g(Bit#(144) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(53, 144, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(53) id, Bit#(144) key);
    actionvalue
      let v <- matchtable_read_ipv6_multicast_route_star_g(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(53) id, Bit#(144) key, Bit#(34) data);
    action
      matchtable_write_ipv6_multicast_route_star_g(key, data);
    endaction
  endfunction

endinstance
interface Ipv6MulticastRouteStarG;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIpv6MulticastRouteStarG  (Ipv6MulticastRouteStarG);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(53, 1024, SizeOf#(Ipv6MulticastRouteStarGReqT), SizeOf#(Ipv6MulticastRouteStarGRspT)) matchTable <- mkMatchTable("ipv6_multicast_route_star_g.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv6_metadata$lkp_ipv6_da = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_da);
    Ipv6MulticastRouteStarGReqT req = Ipv6MulticastRouteStarGReqT {l3_metadata$vrf: l3_metadata$vrf,ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6MulticastRouteStarGRspT resp = unpack(data);
      case (resp._action) matches
        MULTICAST_ROUTE_STAR_G_MISS: begin
          BBRequest req = tagged MulticastRouteStarGMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_ROUTE_SM_STAR_G_HIT: begin
          BBRequest req = tagged MulticastRouteSmStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        MULTICAST_ROUTE_BIDIR_STAR_G_HIT: begin
          BBRequest req = tagged MulticastRouteBidirStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged MulticastRouteStarGMissRspT {pkt: .pkt, l3_metadata$l3_copy: .l3_metadata$l3_copy}: begin
        meta.l3_metadata$l3_copy = tagged Valid l3_metadata$l3_copy;
        MetadataResponse rsp = tagged Ipv6MulticastRouteStarGMulticastRouteStarGMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastRouteSmStarGHitRspT {pkt: .pkt, multicast_metadata$mcast_route_hit: .multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: .multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: .multicast_metadata$mcast_mode}: begin
        meta.multicast_metadata$mcast_route_hit = tagged Valid multicast_metadata$mcast_route_hit;
        meta.multicast_metadata$multicast_route_mc_index = tagged Valid multicast_metadata$multicast_route_mc_index;
        meta.multicast_metadata$mcast_mode = tagged Valid multicast_metadata$mcast_mode;
        MetadataResponse rsp = tagged Ipv6MulticastRouteStarGMulticastRouteSmStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MulticastRouteBidirStarGHitRspT {pkt: .pkt, multicast_metadata$mcast_route_hit: .multicast_metadata$mcast_route_hit, multicast_metadata$multicast_route_mc_index: .multicast_metadata$multicast_route_mc_index, multicast_metadata$mcast_mode: .multicast_metadata$mcast_mode}: begin
        meta.multicast_metadata$mcast_route_hit = tagged Valid multicast_metadata$mcast_route_hit;
        meta.multicast_metadata$multicast_route_mc_index = tagged Valid multicast_metadata$multicast_route_mc_index;
        meta.multicast_metadata$mcast_mode = tagged Valid multicast_metadata$mcast_mode;
        MetadataResponse rsp = tagged Ipv6MulticastRouteStarGMulticastRouteBidirStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== IPV6_RACL ======

typedef struct {
  Bit#(3) padding;
  Bit#(16) acl_metadata$bd_label;
  Bit#(128) ipv6_metadata$lkp_ipv6_sa;
  Bit#(128) ipv6_metadata$lkp_ipv6_da;
  Bit#(8) l3_metadata$lkp_ip_proto;
  Bit#(16) l3_metadata$lkp_l4_sport;
  Bit#(16) l3_metadata$lkp_l4_dport;
} Ipv6RaclReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_RACL,
  NOP,
  RACL_DENY,
  RACL_PERMIT,
  RACL_REDIRECT_NEXTHOP,
  RACL_REDIRECT_ECMP
} Ipv6RaclActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6RaclActionT _action;
  Bit#(14) runtime_acl_stats_index;
  Bit#(1) runtime_acl_copy;
  Bit#(16) runtime_acl_copy_reason;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} Ipv6RaclRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(66)) matchtable_read_ipv6_racl(Bit#(315) msgtype);
import "BDPI" function Action matchtable_write_ipv6_racl(Bit#(315) msgtype, Bit#(66) data);
`endif
instance MatchTableSim#(39, 315, 66);
  function ActionValue#(Bit#(66)) matchtable_read(Bit#(39) id, Bit#(315) key);
    actionvalue
      let v <- matchtable_read_ipv6_racl(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(39) id, Bit#(315) key, Bit#(66) data);
    action
      matchtable_write_ipv6_racl(key, data);
    endaction
  endfunction

endinstance
interface Ipv6Racl;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
endinterface
(* synthesize *)
module mkIpv6Racl  (Ipv6Racl);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(5, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(5, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(39, 512, SizeOf#(Ipv6RaclReqT), SizeOf#(Ipv6RaclRspT)) matchTable <- mkMatchTable("ipv6_racl.dat");
  Vector#(5, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(5) readyChannel = -1;
  for (Integer i=4; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let acl_metadata$bd_label = fromMaybe(?, meta.acl_metadata$bd_label);
    let ipv6_metadata$lkp_ipv6_sa = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_sa);
    let ipv6_metadata$lkp_ipv6_da = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_da);
    let l3_metadata$lkp_ip_proto = fromMaybe(?, meta.l3_metadata$lkp_ip_proto);
    let l3_metadata$lkp_l4_sport = fromMaybe(?, meta.l3_metadata$lkp_l4_sport);
    let l3_metadata$lkp_l4_dport = fromMaybe(?, meta.l3_metadata$lkp_l4_dport);
    Ipv6RaclReqT req = Ipv6RaclReqT {acl_metadata$bd_label: acl_metadata$bd_label,ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa,ipv6_metadata$lkp_ipv6_da: ipv6_metadata$lkp_ipv6_da,l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto,l3_metadata$lkp_l4_sport: l3_metadata$lkp_l4_sport,l3_metadata$lkp_l4_dport: l3_metadata$lkp_l4_dport};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6RaclRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        RACL_DENY: begin
          BBRequest req = tagged RaclDenyReqT {pkt: pkt, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        RACL_PERMIT: begin
          BBRequest req = tagged RaclPermitReqT {pkt: pkt, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        RACL_REDIRECT_NEXTHOP: begin
          BBRequest req = tagged RaclRedirectNexthopReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_nexthop_index: resp.runtime_nexthop_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        RACL_REDIRECT_ECMP: begin
          BBRequest req = tagged RaclRedirectEcmpReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_ecmp_index: resp.runtime_ecmp_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6RaclNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RaclDenyRspT {pkt: .pkt, acl_metadata$racl_deny: .acl_metadata$racl_deny, acl_metadata$acl_copy: .acl_metadata$acl_copy, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index}: begin
        meta.acl_metadata$racl_deny = tagged Valid acl_metadata$racl_deny;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        MetadataResponse rsp = tagged Ipv6RaclRaclDenyRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RaclPermitRspT {pkt: .pkt, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$acl_copy: .acl_metadata$acl_copy, fabric_metadata$reason_code: .fabric_metadata$reason_code}: begin
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        MetadataResponse rsp = tagged Ipv6RaclRaclPermitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RaclRedirectNexthopRspT {pkt: .pkt, acl_metadata$racl_nexthop: .acl_metadata$racl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$racl_redirect: .acl_metadata$racl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$racl_nexthop_type: .acl_metadata$racl_nexthop_type}: begin
        meta.acl_metadata$racl_nexthop = tagged Valid acl_metadata$racl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$racl_redirect = tagged Valid acl_metadata$racl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$racl_nexthop_type = tagged Valid acl_metadata$racl_nexthop_type;
        MetadataResponse rsp = tagged Ipv6RaclRaclRedirectNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RaclRedirectEcmpRspT {pkt: .pkt, acl_metadata$racl_nexthop: .acl_metadata$racl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$racl_redirect: .acl_metadata$racl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$racl_nexthop_type: .acl_metadata$racl_nexthop_type}: begin
        meta.acl_metadata$racl_nexthop = tagged Valid acl_metadata$racl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$racl_redirect = tagged Valid acl_metadata$racl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$racl_nexthop_type = tagged Valid acl_metadata$racl_nexthop_type;
        MetadataResponse rsp = tagged Ipv6RaclRaclRedirectEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
endmodule

// ====== IPV6_SRC_VTEP ======

typedef struct {
  Bit#(4) padding;
  Bit#(16) l3_metadata$vrf;
  Bit#(128) ipv6$srcAddr;
  Bit#(5) tunnel_metadata$ingress_tunnel_type;
} Ipv6SrcVtepReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_SRC_VTEP,
  ON_MISS,
  SRC_VTEP_HIT
} Ipv6SrcVtepActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6SrcVtepActionT _action;
  Bit#(16) runtime_ifindex;
} Ipv6SrcVtepRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv6_src_vtep(Bit#(153) msgtype);
import "BDPI" function Action matchtable_write_ipv6_src_vtep(Bit#(153) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(28, 153, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(28) id, Bit#(153) key);
    actionvalue
      let v <- matchtable_read_ipv6_src_vtep(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(28) id, Bit#(153) key, Bit#(18) data);
    action
      matchtable_write_ipv6_src_vtep(key, data);
    endaction
  endfunction

endinstance
interface Ipv6SrcVtep;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv6SrcVtep  (Ipv6SrcVtep);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(28, 1024, SizeOf#(Ipv6SrcVtepReqT), SizeOf#(Ipv6SrcVtepRspT)) matchTable <- mkMatchTable("ipv6_src_vtep.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv6$srcAddr = fromMaybe(?, meta.ipv6$srcAddr);
    let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
    Ipv6SrcVtepReqT req = Ipv6SrcVtepReqT {l3_metadata$vrf: l3_metadata$vrf,ipv6$srcAddr: ipv6$srcAddr,tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6SrcVtepRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SRC_VTEP_HIT: begin
          BBRequest req = tagged SrcVtepHitReqT {pkt: pkt, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6SrcVtepOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SrcVtepHitRspT {pkt: .pkt, ingress_metadata$ifindex: .ingress_metadata$ifindex}: begin
        meta.ingress_metadata$ifindex = tagged Valid ingress_metadata$ifindex;
        MetadataResponse rsp = tagged Ipv6SrcVtepSrcVtepHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV6_URPF ======

typedef struct {
  Bit#(16) l3_metadata$vrf;
  Bit#(128) ipv6_metadata$lkp_ipv6_sa;
} Ipv6UrpfReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_URPF,
  ON_MISS,
  IPV6_URPF_HIT
} Ipv6UrpfActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6UrpfActionT _action;
  Bit#(16) runtime_urpf_bd_group;
} Ipv6UrpfRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv6_urpf(Bit#(144) msgtype);
import "BDPI" function Action matchtable_write_ipv6_urpf(Bit#(144) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(23, 144, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(23) id, Bit#(144) key);
    actionvalue
      let v <- matchtable_read_ipv6_urpf(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(23) id, Bit#(144) key, Bit#(18) data);
    action
      matchtable_write_ipv6_urpf(key, data);
    endaction
  endfunction

endinstance
interface Ipv6Urpf;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv6Urpf  (Ipv6Urpf);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(23, 1024, SizeOf#(Ipv6UrpfReqT), SizeOf#(Ipv6UrpfRspT)) matchTable <- mkMatchTable("ipv6_urpf.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv6_metadata$lkp_ipv6_sa = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_sa);
    Ipv6UrpfReqT req = Ipv6UrpfReqT {l3_metadata$vrf: l3_metadata$vrf,ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6UrpfRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_URPF_HIT: begin
          BBRequest req = tagged Ipv6UrpfHitReqT {pkt: pkt, ipv6_metadata$ipv6_urpf_mode: ipv6_metadata$ipv6_urpf_mode, runtime_urpf_bd_group: resp.runtime_urpf_bd_group};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged Ipv6UrpfOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6UrpfHitRspT {pkt: .pkt, l3_metadata$urpf_bd_group: .l3_metadata$urpf_bd_group, l3_metadata$urpf_hit: .l3_metadata$urpf_hit, l3_metadata$urpf_mode: .l3_metadata$urpf_mode}: begin
        meta.l3_metadata$urpf_bd_group = tagged Valid l3_metadata$urpf_bd_group;
        meta.l3_metadata$urpf_hit = tagged Valid l3_metadata$urpf_hit;
        meta.l3_metadata$urpf_mode = tagged Valid l3_metadata$urpf_mode;
        MetadataResponse rsp = tagged Ipv6UrpfIpv6UrpfHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== IPV6_URPF_LPM ======

typedef struct {
  Bit#(16) l3_metadata$vrf;
  Bit#(128) ipv6_metadata$lkp_ipv6_sa;
} Ipv6UrpfLpmReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_IPV6_URPF_LPM,
  IPV6_URPF_HIT,
  URPF_MISS
} Ipv6UrpfLpmActionT deriving (Bits, Eq, FShow);
typedef struct {
  Ipv6UrpfLpmActionT _action;
  Bit#(16) runtime_urpf_bd_group;
} Ipv6UrpfLpmRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_ipv6_urpf_lpm(Bit#(144) msgtype);
import "BDPI" function Action matchtable_write_ipv6_urpf_lpm(Bit#(144) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(22, 144, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(22) id, Bit#(144) key);
    actionvalue
      let v <- matchtable_read_ipv6_urpf_lpm(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(22) id, Bit#(144) key, Bit#(18) data);
    action
      matchtable_write_ipv6_urpf_lpm(key, data);
    endaction
  endfunction

endinstance
interface Ipv6UrpfLpm;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIpv6UrpfLpm  (Ipv6UrpfLpm);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(22, 512, SizeOf#(Ipv6UrpfLpmReqT), SizeOf#(Ipv6UrpfLpmRspT)) matchTable <- mkMatchTable("ipv6_urpf_lpm.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$vrf = fromMaybe(?, meta.l3_metadata$vrf);
    let ipv6_metadata$lkp_ipv6_sa = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_sa);
    Ipv6UrpfLpmReqT req = Ipv6UrpfLpmReqT {l3_metadata$vrf: l3_metadata$vrf,ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      Ipv6UrpfLpmRspT resp = unpack(data);
      case (resp._action) matches
        IPV6_URPF_HIT: begin
          BBRequest req = tagged Ipv6UrpfHitReqT {pkt: pkt, ipv6_metadata$ipv6_urpf_mode: ipv6_metadata$ipv6_urpf_mode, runtime_urpf_bd_group: resp.runtime_urpf_bd_group};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        URPF_MISS: begin
          BBRequest req = tagged UrpfMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged Ipv6UrpfHitRspT {pkt: .pkt, l3_metadata$urpf_bd_group: .l3_metadata$urpf_bd_group, l3_metadata$urpf_hit: .l3_metadata$urpf_hit, l3_metadata$urpf_mode: .l3_metadata$urpf_mode}: begin
        meta.l3_metadata$urpf_bd_group = tagged Valid l3_metadata$urpf_bd_group;
        meta.l3_metadata$urpf_hit = tagged Valid l3_metadata$urpf_hit;
        meta.l3_metadata$urpf_mode = tagged Valid l3_metadata$urpf_mode;
        MetadataResponse rsp = tagged Ipv6UrpfLpmIpv6UrpfHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged UrpfMissRspT {pkt: .pkt, l3_metadata$urpf_check_fail: .l3_metadata$urpf_check_fail}: begin
        meta.l3_metadata$urpf_check_fail = tagged Valid l3_metadata$urpf_check_fail;
        MetadataResponse rsp = tagged Ipv6UrpfLpmUrpfMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== LAG_GROUP ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) ingress_metadata$egress_ifindex;
} LagGroupReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_LAG_GROUP,
  SET_LAG_MISS,
  SET_LAG_PORT,
  SET_LAG_REMOTE_PORT
} LagGroupActionT deriving (Bits, Eq, FShow);
typedef struct {
  LagGroupActionT _action;
  Bit#(9) runtime_port;
  Bit#(8) runtime_device;
} LagGroupRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(19)) matchtable_read_lag_group(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_lag_group(Bit#(18) msgtype, Bit#(19) data);
`endif
instance MatchTableSim#(6, 18, 19);
  function ActionValue#(Bit#(19)) matchtable_read(Bit#(6) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_lag_group(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(6) id, Bit#(18) key, Bit#(19) data);
    action
      matchtable_write_lag_group(key, data);
    endaction
  endfunction

endinstance
interface LagGroup;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkLagGroup  (LagGroup);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(6, 1024, SizeOf#(LagGroupReqT), SizeOf#(LagGroupRspT)) matchTable <- mkMatchTable("lag_group.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$egress_ifindex = fromMaybe(?, meta.ingress_metadata$egress_ifindex);
    LagGroupReqT req = LagGroupReqT {ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      LagGroupRspT resp = unpack(data);
      case (resp._action) matches
        SET_LAG_MISS: begin
          BBRequest req = tagged SetLagMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_LAG_PORT: begin
          BBRequest req = tagged SetLagPortReqT {pkt: pkt, runtime_port: resp.runtime_port};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_LAG_REMOTE_PORT: begin
          BBRequest req = tagged SetLagRemotePortReqT {pkt: pkt, runtime_device: resp.runtime_device, runtime_port: resp.runtime_port};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetLagMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged LagGroupSetLagMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetLagPortRspT {pkt: .pkt, standard_metadata$egress_spec: .standard_metadata$egress_spec}: begin
        meta.standard_metadata$egress_spec = tagged Valid standard_metadata$egress_spec;
        MetadataResponse rsp = tagged LagGroupSetLagPortRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetLagRemotePortRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, fabric_metadata$dst_port: .fabric_metadata$dst_port}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.fabric_metadata$dst_port = tagged Valid fabric_metadata$dst_port;
        MetadataResponse rsp = tagged LagGroupSetLagRemotePortRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== LEARN_NOTIFY ======

typedef struct {
  Bit#(7) padding;
  Bit#(1) l2_metadata$l2_src_miss;
  Bit#(16) l2_metadata$l2_src_move;
  Bit#(3) l2_metadata$stp_state;
} LearnNotifyReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_LEARN_NOTIFY,
  NOP,
  GENERATE_LEARN_NOTIFY
} LearnNotifyActionT deriving (Bits, Eq, FShow);
typedef struct {
  LearnNotifyActionT _action;
} LearnNotifyRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_learn_notify(Bit#(27) msgtype);
import "BDPI" function Action matchtable_write_learn_notify(Bit#(27) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(10, 27, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(10) id, Bit#(27) key);
    actionvalue
      let v <- matchtable_read_learn_notify(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(10) id, Bit#(27) key, Bit#(2) data);
    action
      matchtable_write_learn_notify(key, data);
    endaction
  endfunction

endinstance
interface LearnNotify;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkLearnNotify  (LearnNotify);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(10, 512, SizeOf#(LearnNotifyReqT), SizeOf#(LearnNotifyRspT)) matchTable <- mkMatchTable("learn_notify.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l2_metadata$l2_src_miss = fromMaybe(?, meta.l2_metadata$l2_src_miss);
    let l2_metadata$l2_src_move = fromMaybe(?, meta.l2_metadata$l2_src_move);
    let l2_metadata$stp_state = fromMaybe(?, meta.l2_metadata$stp_state);
    LearnNotifyReqT req = LearnNotifyReqT {l2_metadata$l2_src_miss: l2_metadata$l2_src_miss,l2_metadata$l2_src_move: l2_metadata$l2_src_move,l2_metadata$stp_state: l2_metadata$stp_state};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      LearnNotifyRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        GENERATE_LEARN_NOTIFY: begin
          BBRequest req = tagged GenerateLearnNotifyReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged LearnNotifyNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged GenerateLearnNotifyRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged LearnNotifyGenerateLearnNotifyRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== MAC_ACL ======

typedef struct {
  Bit#(16) acl_metadata$if_label;
  Bit#(16) acl_metadata$bd_label;
  Bit#(48) l2_metadata$lkp_mac_sa;
  Bit#(48) l2_metadata$lkp_mac_da;
  Bit#(16) l2_metadata$lkp_mac_type;
} MacAclReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_MAC_ACL,
  NOP,
  ACL_DENY,
  ACL_PERMIT,
  ACL_MIRROR,
  ACL_REDIRECT_NEXTHOP,
  ACL_REDIRECT_ECMP
} MacAclActionT deriving (Bits, Eq, FShow);
typedef struct {
  MacAclActionT _action;
  Bit#(14) runtime_acl_stats_index;
  Bit#(16) runtime_acl_meter_index;
  Bit#(1) runtime_acl_copy;
  Bit#(16) runtime_acl_copy_reason;
  Bit#(32) runtime_session_id;
  Bit#(16) runtime_nexthop_index;
  Bit#(16) runtime_ecmp_index;
} MacAclRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(114)) matchtable_read_mac_acl(Bit#(144) msgtype);
import "BDPI" function Action matchtable_write_mac_acl(Bit#(144) msgtype, Bit#(114) data);
`endif
instance MatchTableSim#(34, 144, 114);
  function ActionValue#(Bit#(114)) matchtable_read(Bit#(34) id, Bit#(144) key);
    actionvalue
      let v <- matchtable_read_mac_acl(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(34) id, Bit#(144) key, Bit#(114) data);
    action
      matchtable_write_mac_acl(key, data);
    endaction
  endfunction

endinstance
interface MacAcl;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
endinterface
(* synthesize *)
module mkMacAcl  (MacAcl);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(6, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(6, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(34, 512, SizeOf#(MacAclReqT), SizeOf#(MacAclRspT)) matchTable <- mkMatchTable("mac_acl.dat");
  Vector#(6, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(6) readyChannel = -1;
  for (Integer i=5; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let acl_metadata$if_label = fromMaybe(?, meta.acl_metadata$if_label);
    let acl_metadata$bd_label = fromMaybe(?, meta.acl_metadata$bd_label);
    let l2_metadata$lkp_mac_sa = fromMaybe(?, meta.l2_metadata$lkp_mac_sa);
    let l2_metadata$lkp_mac_da = fromMaybe(?, meta.l2_metadata$lkp_mac_da);
    let l2_metadata$lkp_mac_type = fromMaybe(?, meta.l2_metadata$lkp_mac_type);
    MacAclReqT req = MacAclReqT {acl_metadata$if_label: acl_metadata$if_label,acl_metadata$bd_label: acl_metadata$bd_label,l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa,l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da,l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      MacAclRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        ACL_DENY: begin
          BBRequest req = tagged AclDenyReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        ACL_PERMIT: begin
          BBRequest req = tagged AclPermitReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_copy: resp.runtime_acl_copy, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        ACL_MIRROR: begin
          BBRequest req = tagged AclMirrorReqT {pkt: pkt, intrinsic_metadata$ingress_global_tstamp: intrinsic_metadata$ingress_global_tstamp, runtime_session_id: resp.runtime_session_id, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        ACL_REDIRECT_NEXTHOP: begin
          BBRequest req = tagged AclRedirectNexthopReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_copy: resp.runtime_acl_copy, runtime_nexthop_index: resp.runtime_nexthop_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        ACL_REDIRECT_ECMP: begin
          BBRequest req = tagged AclRedirectEcmpReqT {pkt: pkt, runtime_acl_copy_reason: resp.runtime_acl_copy_reason, runtime_acl_meter_index: resp.runtime_acl_meter_index, runtime_acl_copy: resp.runtime_acl_copy, runtime_ecmp_index: resp.runtime_ecmp_index, runtime_acl_stats_index: resp.runtime_acl_stats_index};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged MacAclNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclDenyRspT {pkt: .pkt, acl_metadata$acl_deny: .acl_metadata$acl_deny, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_copy: .acl_metadata$acl_copy}: begin
        meta.acl_metadata$acl_deny = tagged Valid acl_metadata$acl_deny;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        MetadataResponse rsp = tagged MacAclAclDenyRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclPermitRspT {pkt: .pkt, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_copy: .acl_metadata$acl_copy}: begin
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        MetadataResponse rsp = tagged MacAclAclPermitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclMirrorRspT {pkt: .pkt, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, meter_metadata$meter_index: .meter_metadata$meter_index, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id}: begin
        meta.i2e_metadata$ingress_tstamp = tagged Valid i2e_metadata$ingress_tstamp;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.i2e_metadata$mirror_session_id = tagged Valid i2e_metadata$mirror_session_id;
        MetadataResponse rsp = tagged MacAclAclMirrorRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclRedirectNexthopRspT {pkt: .pkt, meter_metadata$meter_index: .meter_metadata$meter_index, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$acl_redirect: .acl_metadata$acl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_nexthop: .acl_metadata$acl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_nexthop_type: .acl_metadata$acl_nexthop_type}: begin
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$acl_redirect = tagged Valid acl_metadata$acl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_nexthop = tagged Valid acl_metadata$acl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_nexthop_type = tagged Valid acl_metadata$acl_nexthop_type;
        MetadataResponse rsp = tagged MacAclAclRedirectNexthopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged AclRedirectEcmpRspT {pkt: .pkt, meter_metadata$meter_index: .meter_metadata$meter_index, acl_metadata$acl_stats_index: .acl_metadata$acl_stats_index, acl_metadata$acl_redirect: .acl_metadata$acl_redirect, fabric_metadata$reason_code: .fabric_metadata$reason_code, acl_metadata$acl_nexthop: .acl_metadata$acl_nexthop, acl_metadata$acl_copy: .acl_metadata$acl_copy, acl_metadata$acl_nexthop_type: .acl_metadata$acl_nexthop_type}: begin
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        meta.acl_metadata$acl_stats_index = tagged Valid acl_metadata$acl_stats_index;
        meta.acl_metadata$acl_redirect = tagged Valid acl_metadata$acl_redirect;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.acl_metadata$acl_nexthop = tagged Valid acl_metadata$acl_nexthop;
        meta.acl_metadata$acl_copy = tagged Valid acl_metadata$acl_copy;
        meta.acl_metadata$acl_nexthop_type = tagged Valid acl_metadata$acl_nexthop_type;
        MetadataResponse rsp = tagged MacAclAclRedirectEcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
endmodule

// ====== METER_ACTION ======

typedef struct {
  Bit#(2) meter_metadata$meter_color;
  Bit#(16) meter_metadata$meter_index;
} MeterActionReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_METER_ACTION,
  METER_PERMIT,
  METER_DENY
} MeterActionActionT deriving (Bits, Eq, FShow);
typedef struct {
  MeterActionActionT _action;
} MeterActionRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_meter_action(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_meter_action(Bit#(18) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(74, 18, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(74) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_meter_action(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(74) id, Bit#(18) key, Bit#(2) data);
    action
      matchtable_write_meter_action(key, data);
    endaction
  endfunction

endinstance
interface MeterAction;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkMeterAction  (MeterAction);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(74, 1024, SizeOf#(MeterActionReqT), SizeOf#(MeterActionRspT)) matchTable <- mkMatchTable("meter_action.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let meter_metadata$meter_color = fromMaybe(?, meta.meter_metadata$meter_color);
    let meter_metadata$meter_index = fromMaybe(?, meta.meter_metadata$meter_index);
    MeterActionReqT req = MeterActionReqT {meter_metadata$meter_color: meter_metadata$meter_color,meter_metadata$meter_index: meter_metadata$meter_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      MeterActionRspT resp = unpack(data);
      case (resp._action) matches
        METER_PERMIT: begin
          BBRequest req = tagged MeterPermitReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        METER_DENY: begin
          BBRequest req = tagged MeterDenyReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged MeterPermitRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged MeterActionMeterPermitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MeterDenyRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged MeterActionMeterDenyRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== METER_INDEX ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) meter_metadata$meter_index;
} MeterIndexReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_METER_INDEX,
  NOP
} MeterIndexActionT deriving (Bits, Eq, FShow);
typedef struct {
  MeterIndexActionT _action;
} MeterIndexRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_meter_index(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_meter_index(Bit#(18) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(75, 18, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(75) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_meter_index(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(75) id, Bit#(18) key, Bit#(1) data);
    action
      matchtable_write_meter_index(key, data);
    endaction
  endfunction

endinstance
interface MeterIndex;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkMeterIndex  (MeterIndex);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(75, 1024, SizeOf#(MeterIndexReqT), SizeOf#(MeterIndexRspT)) matchTable <- mkMatchTable("meter_index.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let meter_metadata$meter_index = fromMaybe(?, meta.meter_metadata$meter_index);
    MeterIndexReqT req = MeterIndexReqT {meter_metadata$meter_index: meter_metadata$meter_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      MeterIndexRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged MeterIndexNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== MPLS ======

typedef struct {
  Bit#(5) padding;
  Bit#(20) tunnel_metadata$mpls_label;
  Bit#(Bool) valid_inner_ipv4;
  Bit#(Bool) valid_inner_ipv6;
} MplsReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_MPLS,
  TERMINATE_EOMPLS,
  TERMINATE_VPLS,
  TERMINATE_IPV4_OVER_MPLS,
  TERMINATE_IPV6_OVER_MPLS,
  TERMINATE_PW,
  FORWARD_MPLS
} MplsActionT deriving (Bits, Eq, FShow);
typedef struct {
  MplsActionT _action;
  Bit#(16) runtime_bd;
  Bit#(5) runtime_tunnel_type;
  Bit#(16) runtime_vrf;
  Bit#(16) runtime_ifindex;
  Bit#(16) runtime_nexthop_index;
} MplsRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(72)) matchtable_read_mpls(Bit#(27) msgtype);
import "BDPI" function Action matchtable_write_mpls(Bit#(27) msgtype, Bit#(72) data);
`endif
instance MatchTableSim#(33, 27, 72);
  function ActionValue#(Bit#(72)) matchtable_read(Bit#(33) id, Bit#(27) key);
    actionvalue
      let v <- matchtable_read_mpls(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(33) id, Bit#(27) key, Bit#(72) data);
    action
      matchtable_write_mpls(key, data);
    endaction
  endfunction

endinstance
interface Mpls;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
endinterface
(* synthesize *)
module mkMpls  (Mpls);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(6, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(6, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(33, 1024, SizeOf#(MplsReqT), SizeOf#(MplsRspT)) matchTable <- mkMatchTable("mpls.dat");
  Vector#(6, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(6) readyChannel = -1;
  for (Integer i=5; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$mpls_label = fromMaybe(?, meta.tunnel_metadata$mpls_label);
    let i$n$n$e$r$_$i$p$v$4 = fromMaybe(?, meta.i$n$n$e$r$_$i$p$v$4);
    let i$n$n$e$r$_$i$p$v$6 = fromMaybe(?, meta.i$n$n$e$r$_$i$p$v$6);
    MplsReqT req = MplsReqT {tunnel_metadata$mpls_label: tunnel_metadata$mpls_label,i$n$n$e$r$_$i$p$v$4: i$n$n$e$r$_$i$p$v$4,i$n$n$e$r$_$i$p$v$6: i$n$n$e$r$_$i$p$v$6};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      MplsRspT resp = unpack(data);
      case (resp._action) matches
        TERMINATE_EOMPLS: begin
          BBRequest req = tagged TerminateEomplsReqT {pkt: pkt, inner_ethernet$etherType: inner_ethernet$etherType, runtime_tunnel_type: resp.runtime_tunnel_type, runtime_bd: resp.runtime_bd};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_VPLS: begin
          BBRequest req = tagged TerminateVplsReqT {pkt: pkt, inner_ethernet$etherType: inner_ethernet$etherType, runtime_tunnel_type: resp.runtime_tunnel_type, runtime_bd: resp.runtime_bd};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_IPV4_OVER_MPLS: begin
          BBRequest req = tagged TerminateIpv4OverMplsReqT {pkt: pkt, inner_ipv4$diffserv: inner_ipv4$diffserv, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, inner_ethernet$etherType: inner_ethernet$etherType, inner_ipv4$version: inner_ipv4$version, runtime_tunnel_type: resp.runtime_tunnel_type, runtime_vrf: resp.runtime_vrf};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_IPV6_OVER_MPLS: begin
          BBRequest req = tagged TerminateIpv6OverMplsReqT {pkt: pkt, inner_ipv6$version: inner_ipv6$version, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, inner_ethernet$etherType: inner_ethernet$etherType, inner_ipv6$trafficClass: inner_ipv6$trafficClass, runtime_tunnel_type: resp.runtime_tunnel_type, runtime_vrf: resp.runtime_vrf};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_PW: begin
          BBRequest req = tagged TerminatePwReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        FORWARD_MPLS: begin
          BBRequest req = tagged ForwardMplsReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, runtime_nexthop_index: resp.runtime_nexthop_index};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged TerminateEomplsRspT {pkt: .pkt, tunnel_metadata$ingress_tunnel_type: .tunnel_metadata$ingress_tunnel_type, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type, ingress_metadata$bd: .ingress_metadata$bd}: begin
        meta.tunnel_metadata$ingress_tunnel_type = tagged Valid tunnel_metadata$ingress_tunnel_type;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        meta.ingress_metadata$bd = tagged Valid ingress_metadata$bd;
        MetadataResponse rsp = tagged MplsTerminateEomplsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateVplsRspT {pkt: .pkt, tunnel_metadata$ingress_tunnel_type: .tunnel_metadata$ingress_tunnel_type, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type, ingress_metadata$bd: .ingress_metadata$bd}: begin
        meta.tunnel_metadata$ingress_tunnel_type = tagged Valid tunnel_metadata$ingress_tunnel_type;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        meta.ingress_metadata$bd = tagged Valid ingress_metadata$bd;
        MetadataResponse rsp = tagged MplsTerminateVplsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateIpv4OverMplsRspT {pkt: .pkt, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, tunnel_metadata$ingress_tunnel_type: .tunnel_metadata$ingress_tunnel_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, l3_metadata$vrf: .l3_metadata$vrf, l3_metadata$lkp_ip_version: .l3_metadata$lkp_ip_version, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.tunnel_metadata$ingress_tunnel_type = tagged Valid tunnel_metadata$ingress_tunnel_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        meta.l3_metadata$lkp_ip_tc = tagged Valid l3_metadata$lkp_ip_tc;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.l3_metadata$vrf = tagged Valid l3_metadata$vrf;
        meta.l3_metadata$lkp_ip_version = tagged Valid l3_metadata$lkp_ip_version;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged MplsTerminateIpv4OverMplsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateIpv6OverMplsRspT {pkt: .pkt, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, tunnel_metadata$ingress_tunnel_type: .tunnel_metadata$ingress_tunnel_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, l3_metadata$vrf: .l3_metadata$vrf, l3_metadata$lkp_ip_version: .l3_metadata$lkp_ip_version, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.tunnel_metadata$ingress_tunnel_type = tagged Valid tunnel_metadata$ingress_tunnel_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        meta.l3_metadata$lkp_ip_tc = tagged Valid l3_metadata$lkp_ip_tc;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.l3_metadata$vrf = tagged Valid l3_metadata$vrf;
        meta.l3_metadata$lkp_ip_version = tagged Valid l3_metadata$lkp_ip_version;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged MplsTerminateIpv6OverMplsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminatePwRspT {pkt: .pkt, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged MplsTerminatePwRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged ForwardMplsRspT {pkt: .pkt, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$fib_nexthop: .l3_metadata$fib_nexthop, l3_metadata$fib_hit: .l3_metadata$fib_hit, l3_metadata$fib_nexthop_type: .l3_metadata$fib_nexthop_type, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$fib_nexthop = tagged Valid l3_metadata$fib_nexthop;
        meta.l3_metadata$fib_hit = tagged Valid l3_metadata$fib_hit;
        meta.l3_metadata$fib_nexthop_type = tagged Valid l3_metadata$fib_nexthop_type;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged MplsForwardMplsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
endmodule

// ====== NATIVE_PACKET_OVER_FABRIC ======

typedef struct {
  Bit#(7) padding;
  Bit#(Bool) valid_ipv4;
  Bit#(Bool) valid_ipv6;
} NativePacketOverFabricReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_NATIVE_PACKET_OVER_FABRIC,
  NON_IP_OVER_FABRIC,
  IPV4_OVER_FABRIC,
  IPV6_OVER_FABRIC
} NativePacketOverFabricActionT deriving (Bits, Eq, FShow);
typedef struct {
  NativePacketOverFabricActionT _action;
} NativePacketOverFabricRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_native_packet_over_fabric(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_native_packet_over_fabric(Bit#(9) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(65, 9, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(65) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_native_packet_over_fabric(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(65) id, Bit#(9) key, Bit#(2) data);
    action
      matchtable_write_native_packet_over_fabric(key, data);
    endaction
  endfunction

endinstance
interface NativePacketOverFabric;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkNativePacketOverFabric  (NativePacketOverFabric);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(65, 1024, SizeOf#(NativePacketOverFabricReqT), SizeOf#(NativePacketOverFabricRspT)) matchTable <- mkMatchTable("native_packet_over_fabric.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let i$p$v$6 = fromMaybe(?, meta.i$p$v$6);
    NativePacketOverFabricReqT req = NativePacketOverFabricReqT {i$p$v$4: i$p$v$4,i$p$v$6: i$p$v$6};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      NativePacketOverFabricRspT resp = unpack(data);
      case (resp._action) matches
        NON_IP_OVER_FABRIC: begin
          BBRequest req = tagged NonIpOverFabricReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, ethernet$etherType: ethernet$etherType};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_OVER_FABRIC: begin
          BBRequest req = tagged Ipv4OverFabricReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, ipv4$srcAddr: ipv4$srcAddr, ipv4$dstAddr: ipv4$dstAddr, l3_metadata$lkp_outer_l4_dport: l3_metadata$lkp_outer_l4_dport, ipv4$protocol: ipv4$protocol, l3_metadata$lkp_outer_l4_sport: l3_metadata$lkp_outer_l4_sport};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_OVER_FABRIC: begin
          BBRequest req = tagged Ipv6OverFabricReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, ipv6$srcAddr: ipv6$srcAddr, l3_metadata$lkp_outer_l4_dport: l3_metadata$lkp_outer_l4_dport, ipv6$dstAddr: ipv6$dstAddr, ipv6$nextHdr: ipv6$nextHdr, l3_metadata$lkp_outer_l4_sport: l3_metadata$lkp_outer_l4_sport};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NonIpOverFabricRspT {pkt: .pkt, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged NativePacketOverFabricNonIpOverFabricRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4OverFabricRspT {pkt: .pkt, ipv4_metadata$lkp_ipv4_da: .ipv4_metadata$lkp_ipv4_da, ipv4_metadata$lkp_ipv4_sa: .ipv4_metadata$lkp_ipv4_sa, l3_metadata$lkp_l4_dport: .l3_metadata$lkp_l4_dport, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_sport: .l3_metadata$lkp_l4_sport, l3_metadata$lkp_ip_proto: .l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.ipv4_metadata$lkp_ipv4_da = tagged Valid ipv4_metadata$lkp_ipv4_da;
        meta.ipv4_metadata$lkp_ipv4_sa = tagged Valid ipv4_metadata$lkp_ipv4_sa;
        meta.l3_metadata$lkp_l4_dport = tagged Valid l3_metadata$lkp_l4_dport;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$lkp_l4_sport = tagged Valid l3_metadata$lkp_l4_sport;
        meta.l3_metadata$lkp_ip_proto = tagged Valid l3_metadata$lkp_ip_proto;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged NativePacketOverFabricIpv4OverFabricRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6OverFabricRspT {pkt: .pkt, ipv6_metadata$lkp_ipv6_sa: .ipv6_metadata$lkp_ipv6_sa, ipv6_metadata$lkp_ipv6_da: .ipv6_metadata$lkp_ipv6_da, l3_metadata$lkp_l4_sport: .l3_metadata$lkp_l4_sport, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_dport: .l3_metadata$lkp_l4_dport, l3_metadata$lkp_ip_proto: .l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.ipv6_metadata$lkp_ipv6_sa = tagged Valid ipv6_metadata$lkp_ipv6_sa;
        meta.ipv6_metadata$lkp_ipv6_da = tagged Valid ipv6_metadata$lkp_ipv6_da;
        meta.l3_metadata$lkp_l4_sport = tagged Valid l3_metadata$lkp_l4_sport;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$lkp_l4_dport = tagged Valid l3_metadata$lkp_l4_dport;
        meta.l3_metadata$lkp_ip_proto = tagged Valid l3_metadata$lkp_ip_proto;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged NativePacketOverFabricIpv6OverFabricRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== NEXTHOP ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) l3_metadata$nexthop_index;
} NexthopReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_NEXTHOP,
  NOP,
  SET_NEXTHOP_DETAILS,
  SET_NEXTHOP_DETAILS_FOR_POST_ROUTED_FLOOD
} NexthopActionT deriving (Bits, Eq, FShow);
typedef struct {
  NexthopActionT _action;
  Bit#(16) runtime_ifindex;
  Bit#(16) runtime_bd;
  Bit#(1) runtime_tunnel;
  Bit#(16) runtime_uuc_mc_index;
} NexthopRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(51)) matchtable_read_nexthop(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_nexthop(Bit#(18) msgtype, Bit#(51) data);
`endif
instance MatchTableSim#(58, 18, 51);
  function ActionValue#(Bit#(51)) matchtable_read(Bit#(58) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_nexthop(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(58) id, Bit#(18) key, Bit#(51) data);
    action
      matchtable_write_nexthop(key, data);
    endaction
  endfunction

endinstance
interface Nexthop;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkNexthop  (Nexthop);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(58, 1024, SizeOf#(NexthopReqT), SizeOf#(NexthopRspT)) matchTable <- mkMatchTable("nexthop.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
    NexthopReqT req = NexthopReqT {l3_metadata$nexthop_index: l3_metadata$nexthop_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      NexthopRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_NEXTHOP_DETAILS: begin
          BBRequest req = tagged SetNexthopDetailsReqT {pkt: pkt, runtime_bd: resp.runtime_bd, runtime_tunnel: resp.runtime_tunnel, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_NEXTHOP_DETAILS_FOR_POST_ROUTED_FLOOD: begin
          BBRequest req = tagged SetNexthopDetailsForPostRoutedFloodReqT {pkt: pkt, runtime_uuc_mc_index: resp.runtime_uuc_mc_index, runtime_bd: resp.runtime_bd};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged NexthopNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetNexthopDetailsRspT {pkt: .pkt, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged NexthopSetNexthopDetailsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetNexthopDetailsForPostRoutedFloodRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, ingress_metadata$egress_ifindex: .ingress_metadata$egress_ifindex}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.ingress_metadata$egress_ifindex = tagged Valid ingress_metadata$egress_ifindex;
        MetadataResponse rsp = tagged NexthopSetNexthopDetailsForPostRoutedFloodRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== OUTER_IPV4_MULTICAST ======

typedef struct {
  Bit#(1) multicast_metadata$ipv4_mcast_key_type;
  Bit#(16) multicast_metadata$ipv4_mcast_key;
  Bit#(32) ipv4$srcAddr;
  Bit#(32) ipv4$dstAddr;
} OuterIpv4MulticastReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_OUTER_IPV4_MULTICAST,
  NOP,
  ON_MISS,
  OUTER_MULTICAST_ROUTE_S_G_HIT,
  OUTER_MULTICAST_BRIDGE_S_G_HIT
} OuterIpv4MulticastActionT deriving (Bits, Eq, FShow);
typedef struct {
  OuterIpv4MulticastActionT _action;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_mcast_rpf_group;
} OuterIpv4MulticastRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(35)) matchtable_read_outer_ipv4_multicast(Bit#(81) msgtype);
import "BDPI" function Action matchtable_write_outer_ipv4_multicast(Bit#(81) msgtype, Bit#(35) data);
`endif
instance MatchTableSim#(44, 81, 35);
  function ActionValue#(Bit#(35)) matchtable_read(Bit#(44) id, Bit#(81) key);
    actionvalue
      let v <- matchtable_read_outer_ipv4_multicast(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(44) id, Bit#(81) key, Bit#(35) data);
    action
      matchtable_write_outer_ipv4_multicast(key, data);
    endaction
  endfunction

endinstance
interface OuterIpv4Multicast;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
endinterface
(* synthesize *)
module mkOuterIpv4Multicast  (OuterIpv4Multicast);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(4, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(4, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(44, 1024, SizeOf#(OuterIpv4MulticastReqT), SizeOf#(OuterIpv4MulticastRspT)) matchTable <- mkMatchTable("outer_ipv4_multicast.dat");
  Vector#(4, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(4) readyChannel = -1;
  for (Integer i=3; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let multicast_metadata$ipv4_mcast_key_type = fromMaybe(?, meta.multicast_metadata$ipv4_mcast_key_type);
    let multicast_metadata$ipv4_mcast_key = fromMaybe(?, meta.multicast_metadata$ipv4_mcast_key);
    let ipv4$srcAddr = fromMaybe(?, meta.ipv4$srcAddr);
    let ipv4$dstAddr = fromMaybe(?, meta.ipv4$dstAddr);
    OuterIpv4MulticastReqT req = OuterIpv4MulticastReqT {multicast_metadata$ipv4_mcast_key_type: multicast_metadata$ipv4_mcast_key_type,multicast_metadata$ipv4_mcast_key: multicast_metadata$ipv4_mcast_key,ipv4$srcAddr: ipv4$srcAddr,ipv4$dstAddr: ipv4$dstAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      OuterIpv4MulticastRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_ROUTE_S_G_HIT: begin
          BBRequest req = tagged OuterMulticastRouteSGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_BRIDGE_S_G_HIT: begin
          BBRequest req = tagged OuterMulticastBridgeSGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged OuterIpv4MulticastNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged OuterIpv4MulticastOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastRouteSGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: .multicast_metadata$outer_mcast_route_hit, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.multicast_metadata$outer_mcast_route_hit = tagged Valid multicast_metadata$outer_mcast_route_hit;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv4MulticastOuterMulticastRouteSGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastBridgeSGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv4MulticastOuterMulticastBridgeSGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
endmodule

// ====== OUTER_IPV4_MULTICAST_STAR_G ======

typedef struct {
  Bit#(5) padding;
  Bit#(1) multicast_metadata$ipv4_mcast_key_type;
  Bit#(16) multicast_metadata$ipv4_mcast_key;
  Bit#(32) ipv4$dstAddr;
} OuterIpv4MulticastStarGReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_OUTER_IPV4_MULTICAST_STAR_G,
  NOP,
  OUTER_MULTICAST_ROUTE_SM_STAR_G_HIT,
  OUTER_MULTICAST_ROUTE_BIDIR_STAR_G_HIT,
  OUTER_MULTICAST_BRIDGE_STAR_G_HIT
} OuterIpv4MulticastStarGActionT deriving (Bits, Eq, FShow);
typedef struct {
  OuterIpv4MulticastStarGActionT _action;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_mcast_rpf_group;
} OuterIpv4MulticastStarGRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(35)) matchtable_read_outer_ipv4_multicast_star_g(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_outer_ipv4_multicast_star_g(Bit#(54) msgtype, Bit#(35) data);
`endif
instance MatchTableSim#(43, 54, 35);
  function ActionValue#(Bit#(35)) matchtable_read(Bit#(43) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_outer_ipv4_multicast_star_g(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(43) id, Bit#(54) key, Bit#(35) data);
    action
      matchtable_write_outer_ipv4_multicast_star_g(key, data);
    endaction
  endfunction

endinstance
interface OuterIpv4MulticastStarG;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
endinterface
(* synthesize *)
module mkOuterIpv4MulticastStarG  (OuterIpv4MulticastStarG);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(4, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(4, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(43, 512, SizeOf#(OuterIpv4MulticastStarGReqT), SizeOf#(OuterIpv4MulticastStarGRspT)) matchTable <- mkMatchTable("outer_ipv4_multicast_star_g.dat");
  Vector#(4, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(4) readyChannel = -1;
  for (Integer i=3; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let multicast_metadata$ipv4_mcast_key_type = fromMaybe(?, meta.multicast_metadata$ipv4_mcast_key_type);
    let multicast_metadata$ipv4_mcast_key = fromMaybe(?, meta.multicast_metadata$ipv4_mcast_key);
    let ipv4$dstAddr = fromMaybe(?, meta.ipv4$dstAddr);
    OuterIpv4MulticastStarGReqT req = OuterIpv4MulticastStarGReqT {multicast_metadata$ipv4_mcast_key_type: multicast_metadata$ipv4_mcast_key_type,multicast_metadata$ipv4_mcast_key: multicast_metadata$ipv4_mcast_key,ipv4$dstAddr: ipv4$dstAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      OuterIpv4MulticastStarGRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_ROUTE_SM_STAR_G_HIT: begin
          BBRequest req = tagged OuterMulticastRouteSmStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_ROUTE_BIDIR_STAR_G_HIT: begin
          BBRequest req = tagged OuterMulticastRouteBidirStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_BRIDGE_STAR_G_HIT: begin
          BBRequest req = tagged OuterMulticastBridgeStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged OuterIpv4MulticastStarGNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastRouteSmStarGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: .multicast_metadata$outer_mcast_route_hit, multicast_metadata$outer_mcast_mode: .multicast_metadata$outer_mcast_mode, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.multicast_metadata$outer_mcast_route_hit = tagged Valid multicast_metadata$outer_mcast_route_hit;
        meta.multicast_metadata$outer_mcast_mode = tagged Valid multicast_metadata$outer_mcast_mode;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv4MulticastStarGOuterMulticastRouteSmStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastRouteBidirStarGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: .multicast_metadata$outer_mcast_route_hit, multicast_metadata$outer_mcast_mode: .multicast_metadata$outer_mcast_mode, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.multicast_metadata$outer_mcast_route_hit = tagged Valid multicast_metadata$outer_mcast_route_hit;
        meta.multicast_metadata$outer_mcast_mode = tagged Valid multicast_metadata$outer_mcast_mode;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv4MulticastStarGOuterMulticastRouteBidirStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastBridgeStarGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv4MulticastStarGOuterMulticastBridgeStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
endmodule

// ====== OUTER_IPV6_MULTICAST ======

typedef struct {
  Bit#(6) padding;
  Bit#(1) multicast_metadata$ipv6_mcast_key_type;
  Bit#(16) multicast_metadata$ipv6_mcast_key;
  Bit#(128) ipv6$srcAddr;
  Bit#(128) ipv6$dstAddr;
} OuterIpv6MulticastReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_OUTER_IPV6_MULTICAST,
  NOP,
  ON_MISS,
  OUTER_MULTICAST_ROUTE_S_G_HIT,
  OUTER_MULTICAST_BRIDGE_S_G_HIT
} OuterIpv6MulticastActionT deriving (Bits, Eq, FShow);
typedef struct {
  OuterIpv6MulticastActionT _action;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_mcast_rpf_group;
} OuterIpv6MulticastRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(35)) matchtable_read_outer_ipv6_multicast(Bit#(279) msgtype);
import "BDPI" function Action matchtable_write_outer_ipv6_multicast(Bit#(279) msgtype, Bit#(35) data);
`endif
instance MatchTableSim#(46, 279, 35);
  function ActionValue#(Bit#(35)) matchtable_read(Bit#(46) id, Bit#(279) key);
    actionvalue
      let v <- matchtable_read_outer_ipv6_multicast(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(46) id, Bit#(279) key, Bit#(35) data);
    action
      matchtable_write_outer_ipv6_multicast(key, data);
    endaction
  endfunction

endinstance
interface OuterIpv6Multicast;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
endinterface
(* synthesize *)
module mkOuterIpv6Multicast  (OuterIpv6Multicast);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(4, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(4, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(46, 1024, SizeOf#(OuterIpv6MulticastReqT), SizeOf#(OuterIpv6MulticastRspT)) matchTable <- mkMatchTable("outer_ipv6_multicast.dat");
  Vector#(4, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(4) readyChannel = -1;
  for (Integer i=3; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let multicast_metadata$ipv6_mcast_key_type = fromMaybe(?, meta.multicast_metadata$ipv6_mcast_key_type);
    let multicast_metadata$ipv6_mcast_key = fromMaybe(?, meta.multicast_metadata$ipv6_mcast_key);
    let ipv6$srcAddr = fromMaybe(?, meta.ipv6$srcAddr);
    let ipv6$dstAddr = fromMaybe(?, meta.ipv6$dstAddr);
    OuterIpv6MulticastReqT req = OuterIpv6MulticastReqT {multicast_metadata$ipv6_mcast_key_type: multicast_metadata$ipv6_mcast_key_type,multicast_metadata$ipv6_mcast_key: multicast_metadata$ipv6_mcast_key,ipv6$srcAddr: ipv6$srcAddr,ipv6$dstAddr: ipv6$dstAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      OuterIpv6MulticastRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_ROUTE_S_G_HIT: begin
          BBRequest req = tagged OuterMulticastRouteSGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_BRIDGE_S_G_HIT: begin
          BBRequest req = tagged OuterMulticastBridgeSGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged OuterIpv6MulticastNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged OuterIpv6MulticastOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastRouteSGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: .multicast_metadata$outer_mcast_route_hit, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.multicast_metadata$outer_mcast_route_hit = tagged Valid multicast_metadata$outer_mcast_route_hit;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv6MulticastOuterMulticastRouteSGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastBridgeSGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv6MulticastOuterMulticastBridgeSGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
endmodule

// ====== OUTER_IPV6_MULTICAST_STAR_G ======

typedef struct {
  Bit#(8) padding;
  Bit#(1) multicast_metadata$ipv6_mcast_key_type;
  Bit#(16) multicast_metadata$ipv6_mcast_key;
  Bit#(128) ipv6$dstAddr;
} OuterIpv6MulticastStarGReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_OUTER_IPV6_MULTICAST_STAR_G,
  NOP,
  OUTER_MULTICAST_ROUTE_SM_STAR_G_HIT,
  OUTER_MULTICAST_ROUTE_BIDIR_STAR_G_HIT,
  OUTER_MULTICAST_BRIDGE_STAR_G_HIT
} OuterIpv6MulticastStarGActionT deriving (Bits, Eq, FShow);
typedef struct {
  OuterIpv6MulticastStarGActionT _action;
  Bit#(16) runtime_mc_index;
  Bit#(16) runtime_mcast_rpf_group;
} OuterIpv6MulticastStarGRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(35)) matchtable_read_outer_ipv6_multicast_star_g(Bit#(153) msgtype);
import "BDPI" function Action matchtable_write_outer_ipv6_multicast_star_g(Bit#(153) msgtype, Bit#(35) data);
`endif
instance MatchTableSim#(45, 153, 35);
  function ActionValue#(Bit#(35)) matchtable_read(Bit#(45) id, Bit#(153) key);
    actionvalue
      let v <- matchtable_read_outer_ipv6_multicast_star_g(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(45) id, Bit#(153) key, Bit#(35) data);
    action
      matchtable_write_outer_ipv6_multicast_star_g(key, data);
    endaction
  endfunction

endinstance
interface OuterIpv6MulticastStarG;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
endinterface
(* synthesize *)
module mkOuterIpv6MulticastStarG  (OuterIpv6MulticastStarG);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(4, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(4, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(45, 512, SizeOf#(OuterIpv6MulticastStarGReqT), SizeOf#(OuterIpv6MulticastStarGRspT)) matchTable <- mkMatchTable("outer_ipv6_multicast_star_g.dat");
  Vector#(4, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(4) readyChannel = -1;
  for (Integer i=3; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let multicast_metadata$ipv6_mcast_key_type = fromMaybe(?, meta.multicast_metadata$ipv6_mcast_key_type);
    let multicast_metadata$ipv6_mcast_key = fromMaybe(?, meta.multicast_metadata$ipv6_mcast_key);
    let ipv6$dstAddr = fromMaybe(?, meta.ipv6$dstAddr);
    OuterIpv6MulticastStarGReqT req = OuterIpv6MulticastStarGReqT {multicast_metadata$ipv6_mcast_key_type: multicast_metadata$ipv6_mcast_key_type,multicast_metadata$ipv6_mcast_key: multicast_metadata$ipv6_mcast_key,ipv6$dstAddr: ipv6$dstAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      OuterIpv6MulticastStarGRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_ROUTE_SM_STAR_G_HIT: begin
          BBRequest req = tagged OuterMulticastRouteSmStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_ROUTE_BIDIR_STAR_G_HIT: begin
          BBRequest req = tagged OuterMulticastRouteBidirStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index, runtime_mcast_rpf_group: resp.runtime_mcast_rpf_group};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_MULTICAST_BRIDGE_STAR_G_HIT: begin
          BBRequest req = tagged OuterMulticastBridgeStarGHitReqT {pkt: pkt, runtime_mc_index: resp.runtime_mc_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged OuterIpv6MulticastStarGNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastRouteSmStarGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: .multicast_metadata$outer_mcast_route_hit, multicast_metadata$outer_mcast_mode: .multicast_metadata$outer_mcast_mode, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.multicast_metadata$outer_mcast_route_hit = tagged Valid multicast_metadata$outer_mcast_route_hit;
        meta.multicast_metadata$outer_mcast_mode = tagged Valid multicast_metadata$outer_mcast_mode;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv6MulticastStarGOuterMulticastRouteSmStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastRouteBidirStarGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, multicast_metadata$outer_mcast_route_hit: .multicast_metadata$outer_mcast_route_hit, multicast_metadata$outer_mcast_mode: .multicast_metadata$outer_mcast_mode, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.multicast_metadata$outer_mcast_route_hit = tagged Valid multicast_metadata$outer_mcast_route_hit;
        meta.multicast_metadata$outer_mcast_mode = tagged Valid multicast_metadata$outer_mcast_mode;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv6MulticastStarGOuterMulticastRouteBidirStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterMulticastBridgeStarGHitRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        MetadataResponse rsp = tagged OuterIpv6MulticastStarGOuterMulticastBridgeStarGHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
endmodule

// ====== OUTER_RMAC ======

typedef struct {
  Bit#(5) padding;
  Bit#(10) l3_metadata$rmac_group;
  Bit#(48) ethernet$dstAddr;
} OuterRmacReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_OUTER_RMAC,
  ON_MISS,
  OUTER_RMAC_HIT
} OuterRmacActionT deriving (Bits, Eq, FShow);
typedef struct {
  OuterRmacActionT _action;
} OuterRmacRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_outer_rmac(Bit#(63) msgtype);
import "BDPI" function Action matchtable_write_outer_rmac(Bit#(63) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(24, 63, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(24) id, Bit#(63) key);
    actionvalue
      let v <- matchtable_read_outer_rmac(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(24) id, Bit#(63) key, Bit#(2) data);
    action
      matchtable_write_outer_rmac(key, data);
    endaction
  endfunction

endinstance
interface OuterRmac;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkOuterRmac  (OuterRmac);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(24, 1024, SizeOf#(OuterRmacReqT), SizeOf#(OuterRmacRspT)) matchTable <- mkMatchTable("outer_rmac.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$rmac_group = fromMaybe(?, meta.l3_metadata$rmac_group);
    let ethernet$dstAddr = fromMaybe(?, meta.ethernet$dstAddr);
    OuterRmacReqT req = OuterRmacReqT {l3_metadata$rmac_group: l3_metadata$rmac_group,ethernet$dstAddr: ethernet$dstAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      OuterRmacRspT resp = unpack(data);
      case (resp._action) matches
        ON_MISS: begin
          BBRequest req = tagged OnMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_RMAC_HIT: begin
          BBRequest req = tagged OuterRmacHitReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged OnMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged OuterRmacOnMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterRmacHitRspT {pkt: .pkt, l3_metadata$rmac_hit: .l3_metadata$rmac_hit}: begin
        meta.l3_metadata$rmac_hit = tagged Valid l3_metadata$rmac_hit;
        MetadataResponse rsp = tagged OuterRmacOuterRmacHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== PORT_VLAN_MAPPING ======

typedef struct {
  Bit#(3) padding;
  Bit#(16) ingress_metadata$ifindex;
  Bit#(Bool) valid_vlan_tag_0;
  Bit#(12) vlan_tag_0$vid;
  Bit#(Bool) valid_vlan_tag_1;
  Bit#(12) vlan_tag_1$vid;
} PortVlanMappingReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_PORT_VLAN_MAPPING,
  SET_BD_PROPERTIES,
  PORT_VLAN_MAPPING_MISS
} PortVlanMappingActionT deriving (Bits, Eq, FShow);
typedef struct {
  PortVlanMappingActionT _action;
  Bit#(16) runtime_bd;
  Bit#(16) runtime_vrf;
  Bit#(10) runtime_stp_group;
  Bit#(1) runtime_learning_enabled;
  Bit#(16) runtime_bd_label;
  Bit#(16) runtime_stats_idx;
  Bit#(10) runtime_rmac_group;
  Bit#(1) runtime_ipv4_unicast_enabled;
  Bit#(1) runtime_ipv6_unicast_enabled;
  Bit#(2) runtime_ipv4_urpf_mode;
  Bit#(2) runtime_ipv6_urpf_mode;
  Bit#(1) runtime_igmp_snooping_enabled;
  Bit#(1) runtime_mld_snooping_enabled;
  Bit#(1) runtime_ipv4_multicast_enabled;
  Bit#(1) runtime_ipv6_multicast_enabled;
  Bit#(16) runtime_mrpf_group;
  Bit#(16) runtime_ipv4_mcast_key;
  Bit#(1) runtime_ipv4_mcast_key_type;
  Bit#(16) runtime_ipv6_mcast_key;
  Bit#(1) runtime_ipv6_mcast_key_type;
} PortVlanMappingRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(147)) matchtable_read_port_vlan_mapping(Bit#(45) msgtype);
import "BDPI" function Action matchtable_write_port_vlan_mapping(Bit#(45) msgtype, Bit#(147) data);
`endif
instance MatchTableSim#(4, 45, 147);
  function ActionValue#(Bit#(147)) matchtable_read(Bit#(4) id, Bit#(45) key);
    actionvalue
      let v <- matchtable_read_port_vlan_mapping(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(4) id, Bit#(45) key, Bit#(147) data);
    action
      matchtable_write_port_vlan_mapping(key, data);
    endaction
  endfunction

endinstance
interface PortVlanMapping;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkPortVlanMapping  (PortVlanMapping);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(4, 4096, SizeOf#(PortVlanMappingReqT), SizeOf#(PortVlanMappingRspT)) matchTable <- mkMatchTable("port_vlan_mapping.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$ifindex = fromMaybe(?, meta.ingress_metadata$ifindex);
    let v$l$a$n$_$t$a$g$_$$0$ = fromMaybe(?, meta.v$l$a$n$_$t$a$g$_$$0$);
    let vlan_tag_0$vid = fromMaybe(?, meta.vlan_tag_0$vid);
    let v$l$a$n$_$t$a$g$_$$1$ = fromMaybe(?, meta.v$l$a$n$_$t$a$g$_$$1$);
    let vlan_tag_1$vid = fromMaybe(?, meta.vlan_tag_1$vid);
    PortVlanMappingReqT req = PortVlanMappingReqT {ingress_metadata$ifindex: ingress_metadata$ifindex,v$l$a$n$_$t$a$g$_$$0$: v$l$a$n$_$t$a$g$_$$0$,vlan_tag_0$vid: vlan_tag_0$vid,v$l$a$n$_$t$a$g$_$$1$: v$l$a$n$_$t$a$g$_$$1$,vlan_tag_1$vid: vlan_tag_1$vid};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      PortVlanMappingRspT resp = unpack(data);
      case (resp._action) matches
        SET_BD_PROPERTIES: begin
          BBRequest req = tagged SetBdPropertiesReqT {pkt: pkt, runtime_ipv4_multicast_enabled: resp.runtime_ipv4_multicast_enabled, runtime_igmp_snooping_enabled: resp.runtime_igmp_snooping_enabled, runtime_ipv6_mcast_key: resp.runtime_ipv6_mcast_key, runtime_mrpf_group: resp.runtime_mrpf_group, runtime_ipv4_mcast_key_type: resp.runtime_ipv4_mcast_key_type, runtime_mld_snooping_enabled: resp.runtime_mld_snooping_enabled, runtime_ipv6_multicast_enabled: resp.runtime_ipv6_multicast_enabled, runtime_stats_idx: resp.runtime_stats_idx, runtime_ipv6_urpf_mode: resp.runtime_ipv6_urpf_mode, runtime_ipv4_urpf_mode: resp.runtime_ipv4_urpf_mode, runtime_ipv4_mcast_key: resp.runtime_ipv4_mcast_key, runtime_bd: resp.runtime_bd, runtime_vrf: resp.runtime_vrf, runtime_learning_enabled: resp.runtime_learning_enabled, runtime_ipv6_unicast_enabled: resp.runtime_ipv6_unicast_enabled, runtime_bd_label: resp.runtime_bd_label, runtime_ipv6_mcast_key_type: resp.runtime_ipv6_mcast_key_type, runtime_rmac_group: resp.runtime_rmac_group, runtime_ipv4_unicast_enabled: resp.runtime_ipv4_unicast_enabled, runtime_stp_group: resp.runtime_stp_group};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        PORT_VLAN_MAPPING_MISS: begin
          BBRequest req = tagged PortVlanMappingMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetBdPropertiesRspT {pkt: .pkt, multicast_metadata$ipv4_mcast_key: .multicast_metadata$ipv4_mcast_key, l3_metadata$rmac_group: .l3_metadata$rmac_group, multicast_metadata$igmp_snooping_enabled: .multicast_metadata$igmp_snooping_enabled, multicast_metadata$bd_mrpf_group: .multicast_metadata$bd_mrpf_group, multicast_metadata$ipv4_multicast_enabled: .multicast_metadata$ipv4_multicast_enabled, multicast_metadata$mld_snooping_enabled: .multicast_metadata$mld_snooping_enabled, acl_metadata$bd_label: .acl_metadata$bd_label, l2_metadata$stp_group: .l2_metadata$stp_group, l3_metadata$vrf: .l3_metadata$vrf, ipv6_metadata$ipv6_urpf_mode: .ipv6_metadata$ipv6_urpf_mode, ipv6_metadata$ipv6_unicast_enabled: .ipv6_metadata$ipv6_unicast_enabled, l2_metadata$learning_enabled: .l2_metadata$learning_enabled, ingress_metadata$outer_bd: .ingress_metadata$outer_bd, multicast_metadata$ipv6_mcast_key: .multicast_metadata$ipv6_mcast_key, ingress_metadata$bd: .ingress_metadata$bd, multicast_metadata$ipv4_mcast_key_type: .multicast_metadata$ipv4_mcast_key_type, multicast_metadata$ipv6_mcast_key_type: .multicast_metadata$ipv6_mcast_key_type, ipv4_metadata$ipv4_urpf_mode: .ipv4_metadata$ipv4_urpf_mode, multicast_metadata$ipv6_multicast_enabled: .multicast_metadata$ipv6_multicast_enabled, l2_metadata$bd_stats_idx: .l2_metadata$bd_stats_idx, ipv4_metadata$ipv4_unicast_enabled: .ipv4_metadata$ipv4_unicast_enabled}: begin
        meta.multicast_metadata$ipv4_mcast_key = tagged Valid multicast_metadata$ipv4_mcast_key;
        meta.l3_metadata$rmac_group = tagged Valid l3_metadata$rmac_group;
        meta.multicast_metadata$igmp_snooping_enabled = tagged Valid multicast_metadata$igmp_snooping_enabled;
        meta.multicast_metadata$bd_mrpf_group = tagged Valid multicast_metadata$bd_mrpf_group;
        meta.multicast_metadata$ipv4_multicast_enabled = tagged Valid multicast_metadata$ipv4_multicast_enabled;
        meta.multicast_metadata$mld_snooping_enabled = tagged Valid multicast_metadata$mld_snooping_enabled;
        meta.acl_metadata$bd_label = tagged Valid acl_metadata$bd_label;
        meta.l2_metadata$stp_group = tagged Valid l2_metadata$stp_group;
        meta.l3_metadata$vrf = tagged Valid l3_metadata$vrf;
        meta.ipv6_metadata$ipv6_urpf_mode = tagged Valid ipv6_metadata$ipv6_urpf_mode;
        meta.ipv6_metadata$ipv6_unicast_enabled = tagged Valid ipv6_metadata$ipv6_unicast_enabled;
        meta.l2_metadata$learning_enabled = tagged Valid l2_metadata$learning_enabled;
        meta.ingress_metadata$outer_bd = tagged Valid ingress_metadata$outer_bd;
        meta.multicast_metadata$ipv6_mcast_key = tagged Valid multicast_metadata$ipv6_mcast_key;
        meta.ingress_metadata$bd = tagged Valid ingress_metadata$bd;
        meta.multicast_metadata$ipv4_mcast_key_type = tagged Valid multicast_metadata$ipv4_mcast_key_type;
        meta.multicast_metadata$ipv6_mcast_key_type = tagged Valid multicast_metadata$ipv6_mcast_key_type;
        meta.ipv4_metadata$ipv4_urpf_mode = tagged Valid ipv4_metadata$ipv4_urpf_mode;
        meta.multicast_metadata$ipv6_multicast_enabled = tagged Valid multicast_metadata$ipv6_multicast_enabled;
        meta.l2_metadata$bd_stats_idx = tagged Valid l2_metadata$bd_stats_idx;
        meta.ipv4_metadata$ipv4_unicast_enabled = tagged Valid ipv4_metadata$ipv4_unicast_enabled;
        MetadataResponse rsp = tagged PortVlanMappingSetBdPropertiesRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged PortVlanMappingMissRspT {pkt: .pkt, l2_metadata$port_vlan_mapping_miss: .l2_metadata$port_vlan_mapping_miss}: begin
        meta.l2_metadata$port_vlan_mapping_miss = tagged Valid l2_metadata$port_vlan_mapping_miss;
        MetadataResponse rsp = tagged PortVlanMappingPortVlanMappingMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== QOS ======

typedef struct {
  Bit#(1) padding;
  Bit#(16) acl_metadata$if_label;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
  Bit#(8) l3_metadata$lkp_ip_proto;
  Bit#(8) l3_metadata$lkp_ip_tc;
  Bit#(3) tunnel_metadata$mpls_exp;
  Bit#(8) qos_metadata$outer_dscp;
} QosReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_QOS,
  NOP,
  APPLY_COS_MARKING,
  APPLY_DSCP_MARKING,
  APPLY_TC_MARKING
} QosActionT deriving (Bits, Eq, FShow);
typedef struct {
  QosActionT _action;
  Bit#(3) runtime_cos;
  Bit#(8) runtime_dscp;
  Bit#(3) runtime_tc;
} QosRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(17)) matchtable_read_qos(Bit#(108) msgtype);
import "BDPI" function Action matchtable_write_qos(Bit#(108) msgtype, Bit#(17) data);
`endif
instance MatchTableSim#(37, 108, 17);
  function ActionValue#(Bit#(17)) matchtable_read(Bit#(37) id, Bit#(108) key);
    actionvalue
      let v <- matchtable_read_qos(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(37) id, Bit#(108) key, Bit#(17) data);
    action
      matchtable_write_qos(key, data);
    endaction
  endfunction

endinstance
interface Qos;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
endinterface
(* synthesize *)
module mkQos  (Qos);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(4, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(4, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(37, 512, SizeOf#(QosReqT), SizeOf#(QosRspT)) matchTable <- mkMatchTable("qos.dat");
  Vector#(4, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(4) readyChannel = -1;
  for (Integer i=3; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let acl_metadata$if_label = fromMaybe(?, meta.acl_metadata$if_label);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    let l3_metadata$lkp_ip_proto = fromMaybe(?, meta.l3_metadata$lkp_ip_proto);
    let l3_metadata$lkp_ip_tc = fromMaybe(?, meta.l3_metadata$lkp_ip_tc);
    let tunnel_metadata$mpls_exp = fromMaybe(?, meta.tunnel_metadata$mpls_exp);
    let qos_metadata$outer_dscp = fromMaybe(?, meta.qos_metadata$outer_dscp);
    QosReqT req = QosReqT {acl_metadata$if_label: acl_metadata$if_label,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da,l3_metadata$lkp_ip_proto: l3_metadata$lkp_ip_proto,l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc,tunnel_metadata$mpls_exp: tunnel_metadata$mpls_exp,qos_metadata$outer_dscp: qos_metadata$outer_dscp};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      QosRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        APPLY_COS_MARKING: begin
          BBRequest req = tagged ApplyCosMarkingReqT {pkt: pkt, runtime_cos: resp.runtime_cos};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        APPLY_DSCP_MARKING: begin
          BBRequest req = tagged ApplyDscpMarkingReqT {pkt: pkt, runtime_dscp: resp.runtime_dscp};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        APPLY_TC_MARKING: begin
          BBRequest req = tagged ApplyTcMarkingReqT {pkt: pkt, runtime_tc: resp.runtime_tc};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged QosNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged ApplyCosMarkingRspT {pkt: .pkt, qos_metadata$marked_cos: .qos_metadata$marked_cos}: begin
        meta.qos_metadata$marked_cos = tagged Valid qos_metadata$marked_cos;
        MetadataResponse rsp = tagged QosApplyCosMarkingRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged ApplyDscpMarkingRspT {pkt: .pkt, qos_metadata$marked_dscp: .qos_metadata$marked_dscp}: begin
        meta.qos_metadata$marked_dscp = tagged Valid qos_metadata$marked_dscp;
        MetadataResponse rsp = tagged QosApplyDscpMarkingRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged ApplyTcMarkingRspT {pkt: .pkt, qos_metadata$marked_exp: .qos_metadata$marked_exp}: begin
        meta.qos_metadata$marked_exp = tagged Valid qos_metadata$marked_exp;
        MetadataResponse rsp = tagged QosApplyTcMarkingRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
endmodule

// ====== RMAC ======

typedef struct {
  Bit#(5) padding;
  Bit#(10) l3_metadata$rmac_group;
  Bit#(48) l2_metadata$lkp_mac_da;
} RmacReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_RMAC,
  RMAC_HIT,
  RMAC_MISS
} RmacActionT deriving (Bits, Eq, FShow);
typedef struct {
  RmacActionT _action;
} RmacRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_rmac(Bit#(63) msgtype);
import "BDPI" function Action matchtable_write_rmac(Bit#(63) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(12, 63, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(12) id, Bit#(63) key);
    actionvalue
      let v <- matchtable_read_rmac(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(12) id, Bit#(63) key, Bit#(2) data);
    action
      matchtable_write_rmac(key, data);
    endaction
  endfunction

endinstance
interface Rmac;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkRmac  (Rmac);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(12, 1024, SizeOf#(RmacReqT), SizeOf#(RmacRspT)) matchTable <- mkMatchTable("rmac.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$rmac_group = fromMaybe(?, meta.l3_metadata$rmac_group);
    let l2_metadata$lkp_mac_da = fromMaybe(?, meta.l2_metadata$lkp_mac_da);
    RmacReqT req = RmacReqT {l3_metadata$rmac_group: l3_metadata$rmac_group,l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      RmacRspT resp = unpack(data);
      case (resp._action) matches
        RMAC_HIT: begin
          BBRequest req = tagged RmacHitReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        RMAC_MISS: begin
          BBRequest req = tagged RmacMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged RmacHitRspT {pkt: .pkt, l3_metadata$rmac_hit: .l3_metadata$rmac_hit}: begin
        meta.l3_metadata$rmac_hit = tagged Valid l3_metadata$rmac_hit;
        MetadataResponse rsp = tagged RmacRmacHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RmacMissRspT {pkt: .pkt, l3_metadata$rmac_hit: .l3_metadata$rmac_hit}: begin
        meta.l3_metadata$rmac_hit = tagged Valid l3_metadata$rmac_hit;
        MetadataResponse rsp = tagged RmacRmacMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== SFLOW_ING_TAKE_SAMPLE ======

typedef struct {
  Bit#(6) padding;
  Bit#(32) ingress_metadata$sflow_take_sample;
  Bit#(16) sflow_metadata$sflow_session_id;
} SflowIngTakeSampleReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_SFLOW_ING_TAKE_SAMPLE,
  NOP,
  SFLOW_ING_PKT_TO_CPU
} SflowIngTakeSampleActionT deriving (Bits, Eq, FShow);
typedef struct {
  SflowIngTakeSampleActionT _action;
  Bit#(32) runtime_sflow_i2e_mirror_id;
  Bit#(16) runtime_reason_code;
} SflowIngTakeSampleRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(50)) matchtable_read_sflow_ing_take_sample(Bit#(54) msgtype);
import "BDPI" function Action matchtable_write_sflow_ing_take_sample(Bit#(54) msgtype, Bit#(50) data);
`endif
instance MatchTableSim#(77, 54, 50);
  function ActionValue#(Bit#(50)) matchtable_read(Bit#(77) id, Bit#(54) key);
    actionvalue
      let v <- matchtable_read_sflow_ing_take_sample(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(77) id, Bit#(54) key, Bit#(50) data);
    action
      matchtable_write_sflow_ing_take_sample(key, data);
    endaction
  endfunction

endinstance
interface SflowIngTakeSample;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkSflowIngTakeSample  (SflowIngTakeSample);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(77, 256, SizeOf#(SflowIngTakeSampleReqT), SizeOf#(SflowIngTakeSampleRspT)) matchTable <- mkMatchTable("sflow_ing_take_sample.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$sflow_take_sample = fromMaybe(?, meta.ingress_metadata$sflow_take_sample);
    let sflow_metadata$sflow_session_id = fromMaybe(?, meta.sflow_metadata$sflow_session_id);
    SflowIngTakeSampleReqT req = SflowIngTakeSampleReqT {ingress_metadata$sflow_take_sample: ingress_metadata$sflow_take_sample,sflow_metadata$sflow_session_id: sflow_metadata$sflow_session_id};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      SflowIngTakeSampleRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SFLOW_ING_PKT_TO_CPU: begin
          BBRequest req = tagged SflowIngPktToCpuReqT {pkt: pkt, runtime_sflow_i2e_mirror_id: resp.runtime_sflow_i2e_mirror_id, runtime_reason_code: resp.runtime_reason_code};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SflowIngTakeSampleNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SflowIngPktToCpuRspT {pkt: .pkt, fabric_metadata$reason_code: .fabric_metadata$reason_code, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id}: begin
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        meta.i2e_metadata$mirror_session_id = tagged Valid i2e_metadata$mirror_session_id;
        MetadataResponse rsp = tagged SflowIngTakeSampleSflowIngPktToCpuRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== SFLOW_INGRESS ======

typedef struct {
  Bit#(16) ingress_metadata$ifindex;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
  Bit#(32) ipv4_metadata$lkp_ipv4_da;
  Bit#(Bool) valid_sflow;
} SflowIngressReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_SFLOW_INGRESS,
  NOP,
  SFLOW_ING_SESSION_ENABLE
} SflowIngressActionT deriving (Bits, Eq, FShow);
typedef struct {
  SflowIngressActionT _action;
  Bit#(32) runtime_rate_thr;
  Bit#(16) runtime_session_id;
} SflowIngressRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(50)) matchtable_read_sflow_ingress(Bit#(81) msgtype);
import "BDPI" function Action matchtable_write_sflow_ingress(Bit#(81) msgtype, Bit#(50) data);
`endif
instance MatchTableSim#(76, 81, 50);
  function ActionValue#(Bit#(50)) matchtable_read(Bit#(76) id, Bit#(81) key);
    actionvalue
      let v <- matchtable_read_sflow_ingress(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(76) id, Bit#(81) key, Bit#(50) data);
    action
      matchtable_write_sflow_ingress(key, data);
    endaction
  endfunction

endinstance
interface SflowIngress;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkSflowIngress  (SflowIngress);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(76, 512, SizeOf#(SflowIngressReqT), SizeOf#(SflowIngressRspT)) matchTable <- mkMatchTable("sflow_ingress.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$ifindex = fromMaybe(?, meta.ingress_metadata$ifindex);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    let ipv4_metadata$lkp_ipv4_da = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_da);
    let s$f$l$o$w = fromMaybe(?, meta.s$f$l$o$w);
    SflowIngressReqT req = SflowIngressReqT {ingress_metadata$ifindex: ingress_metadata$ifindex,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa,ipv4_metadata$lkp_ipv4_da: ipv4_metadata$lkp_ipv4_da,s$f$l$o$w: s$f$l$o$w};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      SflowIngressRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SFLOW_ING_SESSION_ENABLE: begin
          BBRequest req = tagged SflowIngSessionEnableReqT {pkt: pkt, runtime_rate_thr: resp.runtime_rate_thr, runtime_session_id: resp.runtime_session_id};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SflowIngressNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SflowIngSessionEnableRspT {pkt: .pkt, sflow_metadata$sflow_session_id: .sflow_metadata$sflow_session_id}: begin
        meta.sflow_metadata$sflow_session_id = tagged Valid sflow_metadata$sflow_session_id;
        MetadataResponse rsp = tagged SflowIngressSflowIngSessionEnableRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== SMAC ======

typedef struct {
  Bit#(8) padding;
  Bit#(16) ingress_metadata$bd;
  Bit#(48) l2_metadata$lkp_mac_sa;
} SmacReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_SMAC,
  NOP,
  SMAC_MISS,
  SMAC_HIT
} SmacActionT deriving (Bits, Eq, FShow);
typedef struct {
  SmacActionT _action;
  Bit#(16) runtime_ifindex;
} SmacRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_smac(Bit#(72) msgtype);
import "BDPI" function Action matchtable_write_smac(Bit#(72) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(8, 72, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(8) id, Bit#(72) key);
    actionvalue
      let v <- matchtable_read_smac(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(8) id, Bit#(72) key, Bit#(18) data);
    action
      matchtable_write_smac(key, data);
    endaction
  endfunction

endinstance
interface Smac;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkSmac  (Smac);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(8, 1024, SizeOf#(SmacReqT), SizeOf#(SmacRspT)) matchTable <- mkMatchTable("smac.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    let l2_metadata$lkp_mac_sa = fromMaybe(?, meta.l2_metadata$lkp_mac_sa);
    SmacReqT req = SmacReqT {ingress_metadata$bd: ingress_metadata$bd,l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      SmacRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SMAC_MISS: begin
          BBRequest req = tagged SmacMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SMAC_HIT: begin
          BBRequest req = tagged SmacHitReqT {pkt: pkt, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SmacNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SmacMissRspT {pkt: .pkt, l2_metadata$l2_src_miss: .l2_metadata$l2_src_miss}: begin
        meta.l2_metadata$l2_src_miss = tagged Valid l2_metadata$l2_src_miss;
        MetadataResponse rsp = tagged SmacSmacMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SmacHitRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SmacSmacHitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== SPANNING_TREE ======

typedef struct {
  Bit#(1) padding;
  Bit#(16) ingress_metadata$ifindex;
  Bit#(10) l2_metadata$stp_group;
} SpanningTreeReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_SPANNING_TREE,
  SET_STP_STATE
} SpanningTreeActionT deriving (Bits, Eq, FShow);
typedef struct {
  SpanningTreeActionT _action;
  Bit#(3) runtime_stp_state;
} SpanningTreeRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(4)) matchtable_read_spanning_tree(Bit#(27) msgtype);
import "BDPI" function Action matchtable_write_spanning_tree(Bit#(27) msgtype, Bit#(4) data);
`endif
instance MatchTableSim#(7, 27, 4);
  function ActionValue#(Bit#(4)) matchtable_read(Bit#(7) id, Bit#(27) key);
    actionvalue
      let v <- matchtable_read_spanning_tree(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(7) id, Bit#(27) key, Bit#(4) data);
    action
      matchtable_write_spanning_tree(key, data);
    endaction
  endfunction

endinstance
interface SpanningTree;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkSpanningTree  (SpanningTree);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(7, 1024, SizeOf#(SpanningTreeReqT), SizeOf#(SpanningTreeRspT)) matchTable <- mkMatchTable("spanning_tree.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ingress_metadata$ifindex = fromMaybe(?, meta.ingress_metadata$ifindex);
    let l2_metadata$stp_group = fromMaybe(?, meta.l2_metadata$stp_group);
    SpanningTreeReqT req = SpanningTreeReqT {ingress_metadata$ifindex: ingress_metadata$ifindex,l2_metadata$stp_group: l2_metadata$stp_group};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      SpanningTreeRspT resp = unpack(data);
      case (resp._action) matches
        SET_STP_STATE: begin
          BBRequest req = tagged SetStpStateReqT {pkt: pkt, runtime_stp_state: resp.runtime_stp_state};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetStpStateRspT {pkt: .pkt, l2_metadata$stp_state: .l2_metadata$stp_state}: begin
        meta.l2_metadata$stp_state = tagged Valid l2_metadata$stp_state;
        MetadataResponse rsp = tagged SpanningTreeSetStpStateRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== STORM_CONTROL ======

typedef struct {
  Bit#(6) padding;
  Bit#(9) standard_metadata$ingress_port;
  Bit#(3) l2_metadata$lkp_pkt_type;
} StormControlReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_STORM_CONTROL,
  NOP,
  SET_STORM_CONTROL_METER
} StormControlActionT deriving (Bits, Eq, FShow);
typedef struct {
  StormControlActionT _action;
  Bit#(32) runtime_meter_idx;
} StormControlRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_storm_control(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_storm_control(Bit#(18) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(60, 18, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(60) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_storm_control(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(60) id, Bit#(18) key, Bit#(34) data);
    action
      matchtable_write_storm_control(key, data);
    endaction
  endfunction

endinstance
interface StormControl;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkStormControl  (StormControl);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(60, 512, SizeOf#(StormControlReqT), SizeOf#(StormControlRspT)) matchTable <- mkMatchTable("storm_control.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let standard_metadata$ingress_port = fromMaybe(?, meta.standard_metadata$ingress_port);
    let l2_metadata$lkp_pkt_type = fromMaybe(?, meta.l2_metadata$lkp_pkt_type);
    StormControlReqT req = StormControlReqT {standard_metadata$ingress_port: standard_metadata$ingress_port,l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      StormControlRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_STORM_CONTROL_METER: begin
          BBRequest req = tagged SetStormControlMeterReqT {pkt: pkt, runtime_meter_idx: resp.runtime_meter_idx};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged StormControlNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetStormControlMeterRspT {pkt: .pkt, meter_metadata$meter_index: .meter_metadata$meter_index}: begin
        meta.meter_metadata$meter_index = tagged Valid meter_metadata$meter_index;
        MetadataResponse rsp = tagged StormControlSetStormControlMeterRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== STORM_CONTROL_STATS ======

typedef struct {
  Bit#(7) padding;
  Bit#(2) meter_metadata$meter_color;
  Bit#(9) standard_metadata$ingress_port;
} StormControlStatsReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_STORM_CONTROL_STATS,
  NOP
} StormControlStatsActionT deriving (Bits, Eq, FShow);
typedef struct {
  StormControlStatsActionT _action;
} StormControlStatsRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_storm_control_stats(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_storm_control_stats(Bit#(18) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(59, 18, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(59) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_storm_control_stats(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(59) id, Bit#(18) key, Bit#(1) data);
    action
      matchtable_write_storm_control_stats(key, data);
    endaction
  endfunction

endinstance
interface StormControlStats;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkStormControlStats  (StormControlStats);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(59, 1024, SizeOf#(StormControlStatsReqT), SizeOf#(StormControlStatsRspT)) matchTable <- mkMatchTable("storm_control_stats.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let meter_metadata$meter_color = fromMaybe(?, meta.meter_metadata$meter_color);
    let standard_metadata$ingress_port = fromMaybe(?, meta.standard_metadata$ingress_port);
    StormControlStatsReqT req = StormControlStatsReqT {meter_metadata$meter_color: meter_metadata$meter_color,standard_metadata$ingress_port: standard_metadata$ingress_port};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      StormControlStatsRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged StormControlStatsNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== SWITCH_CONFIG_PARAMS ======

typedef struct {
} SwitchConfigParamsReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_SWITCH_CONFIG_PARAMS,
  SET_CONFIG_PARAMETERS
} SwitchConfigParamsActionT deriving (Bits, Eq, FShow);
typedef struct {
  SwitchConfigParamsActionT _action;
  Bit#(1) runtime_enable_dod;
} SwitchConfigParamsRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_switch_config_params(Bit#(0) msgtype);
import "BDPI" function Action matchtable_write_switch_config_params(Bit#(0) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(0, 0, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(0) id, Bit#(0) key);
    actionvalue
      let v <- matchtable_read_switch_config_params(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(0) id, Bit#(0) key, Bit#(2) data);
    action
      matchtable_write_switch_config_params(key, data);
    endaction
  endfunction

endinstance
interface SwitchConfigParams;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkSwitchConfigParams  (SwitchConfigParams);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  FIFOF#(MetadataT) metadata_ff <- mkFIFOF;
  rule rl_handle_action_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    packet_ff.enq(pkt);
    metadata_ff.enq(meta);
    let ingress_metadata$ifindex = fromMaybe(?, meta.ingress_metadata$ifindex);
    let intrinsic_metadata$ingress_global_tstamp = fromMaybe(?, meta.intrinsic_metadata$ingress_global_tstamp);
    let standard_metadata$ingress_port = fromMaybe(?, meta.standard_metadata$ingress_port);
    BBRequest req = tagged SetConfigParametersReqT {pkt: pkt, ingress_metadata$ifindex: ingress_metadata$ifindex, intrinsic_metadata$ingress_global_tstamp: intrinsic_metadata$ingress_global_tstamp, standard_metadata$ingress_port: standard_metadata$ingress_port, runtime_enable_dod: resp.runtime_enable_dod};
    bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
  endrule

  rule rl_handle_action_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff).get;
    case (v) matches
      tagged SetConfigParametersRspT {pkt: .pkt, intrinsic_metadata$deflect_on_drop: .intrinsic_metadata$deflect_on_drop, i2e_metadata$ingress_tstamp: .i2e_metadata$ingress_tstamp, ingress_metadata$ingress_port: .ingress_metadata$ingress_port, standard_metadata$egress_spec: .standard_metadata$egress_spec, l2_metadata$same_if_check: .l2_metadata$same_if_check}: begin
        meta.intrinsic_metadata$deflect_on_drop = tagged Valid intrinsic_metadata$deflect_on_drop;
        meta.i2e_metadata$ingress_tstamp = tagged Valid i2e_metadata$ingress_tstamp;
        meta.ingress_metadata$ingress_port = tagged Valid ingress_metadata$ingress_port;
        meta.standard_metadata$egress_spec = tagged Valid standard_metadata$egress_spec;
        meta.l2_metadata$same_if_check = tagged Valid l2_metadata$same_if_check;
        MetadataResponse rsp = tagged SwitchConfigParamsSetConfigParametersRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== SYSTEM_ACL ======

typedef struct {
  Bit#(8) padding;
  Bit#(16) acl_metadata$if_label;
  Bit#(16) acl_metadata$bd_label;
  Bit#(48) l2_metadata$lkp_mac_sa;
  Bit#(48) l2_metadata$lkp_mac_da;
  Bit#(16) l2_metadata$lkp_mac_type;
  Bit#(16) ingress_metadata$ifindex;
  Bit#(1) l2_metadata$port_vlan_mapping_miss;
  Bit#(1) security_metadata$ipsg_check_fail;
  Bit#(1) security_metadata$storm_control_color;
  Bit#(1) acl_metadata$acl_deny;
  Bit#(1) acl_metadata$racl_deny;
  Bit#(1) l3_metadata$urpf_check_fail;
  Bit#(1) ingress_metadata$drop_flag;
  Bit#(1) acl_metadata$acl_copy;
  Bit#(1) l3_metadata$l3_copy;
  Bit#(1) l3_metadata$rmac_hit;
  Bit#(1) l3_metadata$routed;
  Bit#(1) ipv6_metadata$ipv6_src_is_link_local;
  Bit#(16) l2_metadata$same_if_check;
  Bit#(1) tunnel_metadata$tunnel_if_check;
  Bit#(16) l3_metadata$same_bd_check;
  Bit#(8) l3_metadata$lkp_ip_ttl;
  Bit#(3) l2_metadata$stp_state;
  Bit#(1) ingress_metadata$control_frame;
  Bit#(1) ipv4_metadata$ipv4_unicast_enabled;
  Bit#(1) ipv6_metadata$ipv6_unicast_enabled;
  Bit#(16) ingress_metadata$egress_ifindex;
} SystemAclReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_SYSTEM_ACL,
  NOP,
  REDIRECT_TO_CPU,
  COPY_TO_CPU_WITH_REASON,
  COPY_TO_CPU,
  DROP_PACKET,
  DROP_PACKET_WITH_REASON,
  NEGATIVE_MIRROR
} SystemAclActionT deriving (Bits, Eq, FShow);
typedef struct {
  SystemAclActionT _action;
  Bit#(16) runtime_reason_code;
  Bit#(32) runtime_drop_reason;
  Bit#(32) runtime_session_id;
} SystemAclRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(83)) matchtable_read_system_acl(Bit#(243) msgtype);
import "BDPI" function Action matchtable_write_system_acl(Bit#(243) msgtype, Bit#(83) data);
`endif
instance MatchTableSim#(41, 243, 83);
  function ActionValue#(Bit#(83)) matchtable_read(Bit#(41) id, Bit#(243) key);
    actionvalue
      let v <- matchtable_read_system_acl(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(41) id, Bit#(243) key, Bit#(83) data);
    action
      matchtable_write_system_acl(key, data);
    endaction
  endfunction

endinstance
interface SystemAcl;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
endinterface
(* synthesize *)
module mkSystemAcl  (SystemAcl);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(7, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(7, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(41, 512, SizeOf#(SystemAclReqT), SizeOf#(SystemAclRspT)) matchTable <- mkMatchTable("system_acl.dat");
  Vector#(7, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(7) readyChannel = -1;
  for (Integer i=6; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let acl_metadata$if_label = fromMaybe(?, meta.acl_metadata$if_label);
    let acl_metadata$bd_label = fromMaybe(?, meta.acl_metadata$bd_label);
    let l2_metadata$lkp_mac_sa = fromMaybe(?, meta.l2_metadata$lkp_mac_sa);
    let l2_metadata$lkp_mac_da = fromMaybe(?, meta.l2_metadata$lkp_mac_da);
    let l2_metadata$lkp_mac_type = fromMaybe(?, meta.l2_metadata$lkp_mac_type);
    let ingress_metadata$ifindex = fromMaybe(?, meta.ingress_metadata$ifindex);
    let l2_metadata$port_vlan_mapping_miss = fromMaybe(?, meta.l2_metadata$port_vlan_mapping_miss);
    let security_metadata$ipsg_check_fail = fromMaybe(?, meta.security_metadata$ipsg_check_fail);
    let security_metadata$storm_control_color = fromMaybe(?, meta.security_metadata$storm_control_color);
    let acl_metadata$acl_deny = fromMaybe(?, meta.acl_metadata$acl_deny);
    let acl_metadata$racl_deny = fromMaybe(?, meta.acl_metadata$racl_deny);
    let l3_metadata$urpf_check_fail = fromMaybe(?, meta.l3_metadata$urpf_check_fail);
    let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
    let acl_metadata$acl_copy = fromMaybe(?, meta.acl_metadata$acl_copy);
    let l3_metadata$l3_copy = fromMaybe(?, meta.l3_metadata$l3_copy);
    let l3_metadata$rmac_hit = fromMaybe(?, meta.l3_metadata$rmac_hit);
    let l3_metadata$routed = fromMaybe(?, meta.l3_metadata$routed);
    let ipv6_metadata$ipv6_src_is_link_local = fromMaybe(?, meta.ipv6_metadata$ipv6_src_is_link_local);
    let l2_metadata$same_if_check = fromMaybe(?, meta.l2_metadata$same_if_check);
    let tunnel_metadata$tunnel_if_check = fromMaybe(?, meta.tunnel_metadata$tunnel_if_check);
    let l3_metadata$same_bd_check = fromMaybe(?, meta.l3_metadata$same_bd_check);
    let l3_metadata$lkp_ip_ttl = fromMaybe(?, meta.l3_metadata$lkp_ip_ttl);
    let l2_metadata$stp_state = fromMaybe(?, meta.l2_metadata$stp_state);
    let ingress_metadata$control_frame = fromMaybe(?, meta.ingress_metadata$control_frame);
    let ipv4_metadata$ipv4_unicast_enabled = fromMaybe(?, meta.ipv4_metadata$ipv4_unicast_enabled);
    let ipv6_metadata$ipv6_unicast_enabled = fromMaybe(?, meta.ipv6_metadata$ipv6_unicast_enabled);
    let ingress_metadata$egress_ifindex = fromMaybe(?, meta.ingress_metadata$egress_ifindex);
    SystemAclReqT req = SystemAclReqT {acl_metadata$if_label: acl_metadata$if_label,acl_metadata$bd_label: acl_metadata$bd_label,l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa,l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da,l2_metadata$lkp_mac_type: l2_metadata$lkp_mac_type,ingress_metadata$ifindex: ingress_metadata$ifindex,l2_metadata$port_vlan_mapping_miss: l2_metadata$port_vlan_mapping_miss,security_metadata$ipsg_check_fail: security_metadata$ipsg_check_fail,security_metadata$storm_control_color: security_metadata$storm_control_color,acl_metadata$acl_deny: acl_metadata$acl_deny,acl_metadata$racl_deny: acl_metadata$racl_deny,l3_metadata$urpf_check_fail: l3_metadata$urpf_check_fail,ingress_metadata$drop_flag: ingress_metadata$drop_flag,acl_metadata$acl_copy: acl_metadata$acl_copy,l3_metadata$l3_copy: l3_metadata$l3_copy,l3_metadata$rmac_hit: l3_metadata$rmac_hit,l3_metadata$routed: l3_metadata$routed,ipv6_metadata$ipv6_src_is_link_local: ipv6_metadata$ipv6_src_is_link_local,l2_metadata$same_if_check: l2_metadata$same_if_check,tunnel_metadata$tunnel_if_check: tunnel_metadata$tunnel_if_check,l3_metadata$same_bd_check: l3_metadata$same_bd_check,l3_metadata$lkp_ip_ttl: l3_metadata$lkp_ip_ttl,l2_metadata$stp_state: l2_metadata$stp_state,ingress_metadata$control_frame: ingress_metadata$control_frame,ipv4_metadata$ipv4_unicast_enabled: ipv4_metadata$ipv4_unicast_enabled,ipv6_metadata$ipv6_unicast_enabled: ipv6_metadata$ipv6_unicast_enabled,ingress_metadata$egress_ifindex: ingress_metadata$egress_ifindex};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      SystemAclRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        REDIRECT_TO_CPU: begin
          BBRequest req = tagged RedirectToCpuReqT {pkt: pkt, runtime_reason_code: resp.runtime_reason_code};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        COPY_TO_CPU_WITH_REASON: begin
          BBRequest req = tagged CopyToCpuWithReasonReqT {pkt: pkt, runtime_reason_code: resp.runtime_reason_code};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        COPY_TO_CPU: begin
          BBRequest req = tagged CopyToCpuReqT {pkt: pkt};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        DROP_PACKET: begin
          BBRequest req = tagged DropPacketReqT {pkt: pkt};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        DROP_PACKET_WITH_REASON: begin
          BBRequest req = tagged DropPacketWithReasonReqT {pkt: pkt, runtime_drop_reason: resp.runtime_drop_reason};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        NEGATIVE_MIRROR: begin
          BBRequest req = tagged NegativeMirrorReqT {pkt: pkt, runtime_session_id: resp.runtime_session_id};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SystemAclNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RedirectToCpuRspT {pkt: .pkt, fabric_metadata$dst_device: .fabric_metadata$dst_device, fabric_metadata$reason_code: .fabric_metadata$reason_code}: begin
        meta.fabric_metadata$dst_device = tagged Valid fabric_metadata$dst_device;
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        MetadataResponse rsp = tagged SystemAclRedirectToCpuRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged CopyToCpuWithReasonRspT {pkt: .pkt, fabric_metadata$reason_code: .fabric_metadata$reason_code}: begin
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        MetadataResponse rsp = tagged SystemAclCopyToCpuWithReasonRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged CopyToCpuRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SystemAclCopyToCpuRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DropPacketRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SystemAclDropPacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DropPacketWithReasonRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SystemAclDropPacketWithReasonRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged NegativeMirrorRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged SystemAclNegativeMirrorRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
endmodule

// ====== TUNNEL ======

typedef struct {
  Bit#(5) padding;
  Bit#(24) tunnel_metadata$tunnel_vni;
  Bit#(5) tunnel_metadata$ingress_tunnel_type;
  Bit#(Bool) valid_inner_ipv4;
  Bit#(Bool) valid_inner_ipv6;
} TunnelReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL,
  NOP,
  TUNNEL_LOOKUP_MISS,
  TERMINATE_TUNNEL_INNER_NON_IP,
  TERMINATE_TUNNEL_INNER_ETHERNET_IPV4,
  TERMINATE_TUNNEL_INNER_IPV4,
  TERMINATE_TUNNEL_INNER_ETHERNET_IPV6,
  TERMINATE_TUNNEL_INNER_IPV6
} TunnelActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelActionT _action;
  Bit#(16) runtime_bd;
  Bit#(16) runtime_bd_label;
  Bit#(16) runtime_stats_idx;
  Bit#(16) runtime_vrf;
  Bit#(10) runtime_rmac_group;
  Bit#(1) runtime_ipv4_unicast_enabled;
  Bit#(2) runtime_ipv4_urpf_mode;
  Bit#(1) runtime_igmp_snooping_enabled;
  Bit#(1) runtime_ipv4_multicast_enabled;
  Bit#(16) runtime_mrpf_group;
  Bit#(1) runtime_ipv6_unicast_enabled;
  Bit#(2) runtime_ipv6_urpf_mode;
  Bit#(1) runtime_mld_snooping_enabled;
  Bit#(1) runtime_ipv6_multicast_enabled;
} TunnelRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(103)) matchtable_read_tunnel(Bit#(36) msgtype);
import "BDPI" function Action matchtable_write_tunnel(Bit#(36) msgtype, Bit#(103) data);
`endif
instance MatchTableSim#(29, 36, 103);
  function ActionValue#(Bit#(103)) matchtable_read(Bit#(29) id, Bit#(36) key);
    actionvalue
      let v <- matchtable_read_tunnel(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(29) id, Bit#(36) key, Bit#(103) data);
    action
      matchtable_write_tunnel(key, data);
    endaction
  endfunction

endinstance
interface Tunnel;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
endinterface
(* synthesize *)
module mkTunnel  (Tunnel);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(7, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(7, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(29, 1024, SizeOf#(TunnelReqT), SizeOf#(TunnelRspT)) matchTable <- mkMatchTable("tunnel.dat");
  Vector#(7, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(7) readyChannel = -1;
  for (Integer i=6; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$tunnel_vni = fromMaybe(?, meta.tunnel_metadata$tunnel_vni);
    let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
    let i$n$n$e$r$_$i$p$v$4 = fromMaybe(?, meta.i$n$n$e$r$_$i$p$v$4);
    let i$n$n$e$r$_$i$p$v$6 = fromMaybe(?, meta.i$n$n$e$r$_$i$p$v$6);
    TunnelReqT req = TunnelReqT {tunnel_metadata$tunnel_vni: tunnel_metadata$tunnel_vni,tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type,i$n$n$e$r$_$i$p$v$4: i$n$n$e$r$_$i$p$v$4,i$n$n$e$r$_$i$p$v$6: i$n$n$e$r$_$i$p$v$6};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        TUNNEL_LOOKUP_MISS: begin
          BBRequest req = tagged TunnelLookupMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_TUNNEL_INNER_NON_IP: begin
          BBRequest req = tagged TerminateTunnelInnerNonIpReqT {pkt: pkt, inner_ethernet$etherType: inner_ethernet$etherType, runtime_bd_label: resp.runtime_bd_label, runtime_bd: resp.runtime_bd, runtime_stats_idx: resp.runtime_stats_idx};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_TUNNEL_INNER_ETHERNET_IPV4: begin
          BBRequest req = tagged TerminateTunnelInnerEthernetIpv4ReqT {pkt: pkt, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, inner_ipv4$version: inner_ipv4$version, inner_ethernet$etherType: inner_ethernet$etherType, inner_ipv4$diffserv: inner_ipv4$diffserv, runtime_ipv4_multicast_enabled: resp.runtime_ipv4_multicast_enabled, runtime_igmp_snooping_enabled: resp.runtime_igmp_snooping_enabled, runtime_mrpf_group: resp.runtime_mrpf_group, runtime_stats_idx: resp.runtime_stats_idx, runtime_ipv4_urpf_mode: resp.runtime_ipv4_urpf_mode, runtime_bd: resp.runtime_bd, runtime_vrf: resp.runtime_vrf, runtime_bd_label: resp.runtime_bd_label, runtime_rmac_group: resp.runtime_rmac_group, runtime_ipv4_unicast_enabled: resp.runtime_ipv4_unicast_enabled};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_TUNNEL_INNER_IPV4: begin
          BBRequest req = tagged TerminateTunnelInnerIpv4ReqT {pkt: pkt, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, inner_ipv4$diffserv: inner_ipv4$diffserv, inner_ipv4$version: inner_ipv4$version, runtime_ipv4_multicast_enabled: resp.runtime_ipv4_multicast_enabled, runtime_mrpf_group: resp.runtime_mrpf_group, runtime_ipv4_urpf_mode: resp.runtime_ipv4_urpf_mode, runtime_vrf: resp.runtime_vrf, runtime_rmac_group: resp.runtime_rmac_group, runtime_ipv4_unicast_enabled: resp.runtime_ipv4_unicast_enabled};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_TUNNEL_INNER_ETHERNET_IPV6: begin
          BBRequest req = tagged TerminateTunnelInnerEthernetIpv6ReqT {pkt: pkt, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, inner_ipv6$trafficClass: inner_ipv6$trafficClass, inner_ethernet$etherType: inner_ethernet$etherType, inner_ipv6$version: inner_ipv6$version, runtime_mrpf_group: resp.runtime_mrpf_group, runtime_mld_snooping_enabled: resp.runtime_mld_snooping_enabled, runtime_ipv6_multicast_enabled: resp.runtime_ipv6_multicast_enabled, runtime_stats_idx: resp.runtime_stats_idx, runtime_ipv6_urpf_mode: resp.runtime_ipv6_urpf_mode, runtime_bd: resp.runtime_bd, runtime_vrf: resp.runtime_vrf, runtime_ipv6_unicast_enabled: resp.runtime_ipv6_unicast_enabled, runtime_bd_label: resp.runtime_bd_label, runtime_rmac_group: resp.runtime_rmac_group};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        TERMINATE_TUNNEL_INNER_IPV6: begin
          BBRequest req = tagged TerminateTunnelInnerIpv6ReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, inner_ipv6$dstAddr: inner_ipv6$dstAddr, inner_ipv6$srcAddr: inner_ipv6$srcAddr, l3_metadata$lkp_ip_tc: l3_metadata$lkp_ip_tc, inner_ipv6$trafficClass: inner_ipv6$trafficClass, inner_ipv6$version: inner_ipv6$version, runtime_mrpf_group: resp.runtime_mrpf_group, runtime_ipv6_multicast_enabled: resp.runtime_ipv6_multicast_enabled, runtime_ipv6_urpf_mode: resp.runtime_ipv6_urpf_mode, runtime_vrf: resp.runtime_vrf, runtime_ipv6_unicast_enabled: resp.runtime_ipv6_unicast_enabled, runtime_rmac_group: resp.runtime_rmac_group};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TunnelLookupMissRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelTunnelLookupMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateTunnelInnerNonIpRspT {pkt: .pkt, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, ingress_metadata$bd: .ingress_metadata$bd, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type, acl_metadata$bd_label: .acl_metadata$bd_label, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, l2_metadata$bd_stats_idx: .l2_metadata$bd_stats_idx}: begin
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.ingress_metadata$bd = tagged Valid ingress_metadata$bd;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        meta.acl_metadata$bd_label = tagged Valid acl_metadata$bd_label;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.l2_metadata$bd_stats_idx = tagged Valid l2_metadata$bd_stats_idx;
        MetadataResponse rsp = tagged TunnelTerminateTunnelInnerNonIpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateTunnelInnerEthernetIpv4RspT {pkt: .pkt, l3_metadata$rmac_group: .l3_metadata$rmac_group, multicast_metadata$igmp_snooping_enabled: .multicast_metadata$igmp_snooping_enabled, multicast_metadata$bd_mrpf_group: .multicast_metadata$bd_mrpf_group, multicast_metadata$ipv4_multicast_enabled: .multicast_metadata$ipv4_multicast_enabled, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type, acl_metadata$bd_label: .acl_metadata$bd_label, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, l3_metadata$vrf: .l3_metadata$vrf, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, l3_metadata$lkp_ip_version: .l3_metadata$lkp_ip_version, qos_metadata$outer_dscp: .qos_metadata$outer_dscp, ingress_metadata$bd: .ingress_metadata$bd, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, ipv4_metadata$ipv4_urpf_mode: .ipv4_metadata$ipv4_urpf_mode, l2_metadata$bd_stats_idx: .l2_metadata$bd_stats_idx, ipv4_metadata$ipv4_unicast_enabled: .ipv4_metadata$ipv4_unicast_enabled}: begin
        meta.l3_metadata$rmac_group = tagged Valid l3_metadata$rmac_group;
        meta.multicast_metadata$igmp_snooping_enabled = tagged Valid multicast_metadata$igmp_snooping_enabled;
        meta.multicast_metadata$bd_mrpf_group = tagged Valid multicast_metadata$bd_mrpf_group;
        meta.multicast_metadata$ipv4_multicast_enabled = tagged Valid multicast_metadata$ipv4_multicast_enabled;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        meta.acl_metadata$bd_label = tagged Valid acl_metadata$bd_label;
        meta.l3_metadata$lkp_ip_tc = tagged Valid l3_metadata$lkp_ip_tc;
        meta.l3_metadata$vrf = tagged Valid l3_metadata$vrf;
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.l3_metadata$lkp_ip_version = tagged Valid l3_metadata$lkp_ip_version;
        meta.qos_metadata$outer_dscp = tagged Valid qos_metadata$outer_dscp;
        meta.ingress_metadata$bd = tagged Valid ingress_metadata$bd;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.ipv4_metadata$ipv4_urpf_mode = tagged Valid ipv4_metadata$ipv4_urpf_mode;
        meta.l2_metadata$bd_stats_idx = tagged Valid l2_metadata$bd_stats_idx;
        meta.ipv4_metadata$ipv4_unicast_enabled = tagged Valid ipv4_metadata$ipv4_unicast_enabled;
        MetadataResponse rsp = tagged TunnelTerminateTunnelInnerEthernetIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateTunnelInnerIpv4RspT {pkt: .pkt, l3_metadata$rmac_group: .l3_metadata$rmac_group, ipv4_metadata$ipv4_urpf_mode: .ipv4_metadata$ipv4_urpf_mode, multicast_metadata$bd_mrpf_group: .multicast_metadata$bd_mrpf_group, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, l3_metadata$vrf: .l3_metadata$vrf, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, multicast_metadata$ipv4_multicast_enabled: .multicast_metadata$ipv4_multicast_enabled, qos_metadata$outer_dscp: .qos_metadata$outer_dscp, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, ipv4_metadata$ipv4_unicast_enabled: .ipv4_metadata$ipv4_unicast_enabled, l3_metadata$lkp_ip_version: .l3_metadata$lkp_ip_version, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l3_metadata$rmac_group = tagged Valid l3_metadata$rmac_group;
        meta.ipv4_metadata$ipv4_urpf_mode = tagged Valid ipv4_metadata$ipv4_urpf_mode;
        meta.multicast_metadata$bd_mrpf_group = tagged Valid multicast_metadata$bd_mrpf_group;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$lkp_ip_tc = tagged Valid l3_metadata$lkp_ip_tc;
        meta.l3_metadata$vrf = tagged Valid l3_metadata$vrf;
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.multicast_metadata$ipv4_multicast_enabled = tagged Valid multicast_metadata$ipv4_multicast_enabled;
        meta.qos_metadata$outer_dscp = tagged Valid qos_metadata$outer_dscp;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.ipv4_metadata$ipv4_unicast_enabled = tagged Valid ipv4_metadata$ipv4_unicast_enabled;
        meta.l3_metadata$lkp_ip_version = tagged Valid l3_metadata$lkp_ip_version;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged TunnelTerminateTunnelInnerIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateTunnelInnerEthernetIpv6RspT {pkt: .pkt, l3_metadata$rmac_group: .l3_metadata$rmac_group, multicast_metadata$bd_mrpf_group: .multicast_metadata$bd_mrpf_group, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type, acl_metadata$bd_label: .acl_metadata$bd_label, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, l3_metadata$vrf: .l3_metadata$vrf, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, ipv6_metadata$ipv6_unicast_enabled: .ipv6_metadata$ipv6_unicast_enabled, ipv6_metadata$ipv6_urpf_mode: .ipv6_metadata$ipv6_urpf_mode, qos_metadata$outer_dscp: .qos_metadata$outer_dscp, ingress_metadata$bd: .ingress_metadata$bd, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, multicast_metadata$ipv6_multicast_enabled: .multicast_metadata$ipv6_multicast_enabled, l2_metadata$bd_stats_idx: .l2_metadata$bd_stats_idx, l3_metadata$lkp_ip_version: .l3_metadata$lkp_ip_version, multicast_metadata$mld_snooping_enabled: .multicast_metadata$mld_snooping_enabled}: begin
        meta.l3_metadata$rmac_group = tagged Valid l3_metadata$rmac_group;
        meta.multicast_metadata$bd_mrpf_group = tagged Valid multicast_metadata$bd_mrpf_group;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        meta.acl_metadata$bd_label = tagged Valid acl_metadata$bd_label;
        meta.l3_metadata$lkp_ip_tc = tagged Valid l3_metadata$lkp_ip_tc;
        meta.l3_metadata$vrf = tagged Valid l3_metadata$vrf;
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.ipv6_metadata$ipv6_unicast_enabled = tagged Valid ipv6_metadata$ipv6_unicast_enabled;
        meta.ipv6_metadata$ipv6_urpf_mode = tagged Valid ipv6_metadata$ipv6_urpf_mode;
        meta.qos_metadata$outer_dscp = tagged Valid qos_metadata$outer_dscp;
        meta.ingress_metadata$bd = tagged Valid ingress_metadata$bd;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.multicast_metadata$ipv6_multicast_enabled = tagged Valid multicast_metadata$ipv6_multicast_enabled;
        meta.l2_metadata$bd_stats_idx = tagged Valid l2_metadata$bd_stats_idx;
        meta.l3_metadata$lkp_ip_version = tagged Valid l3_metadata$lkp_ip_version;
        meta.multicast_metadata$mld_snooping_enabled = tagged Valid multicast_metadata$mld_snooping_enabled;
        MetadataResponse rsp = tagged TunnelTerminateTunnelInnerEthernetIpv6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TerminateTunnelInnerIpv6RspT {pkt: .pkt, l3_metadata$rmac_group: .l3_metadata$rmac_group, qos_metadata$outer_dscp: .qos_metadata$outer_dscp, multicast_metadata$bd_mrpf_group: .multicast_metadata$bd_mrpf_group, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, l3_metadata$vrf: .l3_metadata$vrf, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, ipv6_metadata$ipv6_unicast_enabled: .ipv6_metadata$ipv6_unicast_enabled, ipv6_metadata$lkp_ipv6_sa: .ipv6_metadata$lkp_ipv6_sa, ipv6_metadata$ipv6_urpf_mode: .ipv6_metadata$ipv6_urpf_mode, ipv6_metadata$lkp_ipv6_da: .ipv6_metadata$lkp_ipv6_da, tunnel_metadata$tunnel_terminate: .tunnel_metadata$tunnel_terminate, multicast_metadata$ipv6_multicast_enabled: .multicast_metadata$ipv6_multicast_enabled, l3_metadata$lkp_ip_version: .l3_metadata$lkp_ip_version, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l3_metadata$rmac_group = tagged Valid l3_metadata$rmac_group;
        meta.qos_metadata$outer_dscp = tagged Valid qos_metadata$outer_dscp;
        meta.multicast_metadata$bd_mrpf_group = tagged Valid multicast_metadata$bd_mrpf_group;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$lkp_ip_tc = tagged Valid l3_metadata$lkp_ip_tc;
        meta.l3_metadata$vrf = tagged Valid l3_metadata$vrf;
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.ipv6_metadata$ipv6_unicast_enabled = tagged Valid ipv6_metadata$ipv6_unicast_enabled;
        meta.ipv6_metadata$lkp_ipv6_sa = tagged Valid ipv6_metadata$lkp_ipv6_sa;
        meta.ipv6_metadata$ipv6_urpf_mode = tagged Valid ipv6_metadata$ipv6_urpf_mode;
        meta.ipv6_metadata$lkp_ipv6_da = tagged Valid ipv6_metadata$lkp_ipv6_da;
        meta.tunnel_metadata$tunnel_terminate = tagged Valid tunnel_metadata$tunnel_terminate;
        meta.multicast_metadata$ipv6_multicast_enabled = tagged Valid multicast_metadata$ipv6_multicast_enabled;
        meta.l3_metadata$lkp_ip_version = tagged Valid l3_metadata$lkp_ip_version;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged TunnelTerminateTunnelInnerIpv6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
endmodule

// ====== TUNNEL_LOOKUP_MISS ======

typedef struct {
  Bit#(7) padding;
  Bit#(Bool) valid_ipv4;
  Bit#(Bool) valid_ipv6;
} TunnelLookupMissReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_LOOKUP_MISS,
  NON_IP_TUNNEL_LOOKUP_MISS,
  IPV4_TUNNEL_LOOKUP_MISS,
  IPV6_TUNNEL_LOOKUP_MISS
} TunnelLookupMissActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelLookupMissActionT _action;
} TunnelLookupMissRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_tunnel_lookup_miss(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_tunnel_lookup_miss(Bit#(9) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(31, 9, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(31) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_tunnel_lookup_miss(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(31) id, Bit#(9) key, Bit#(2) data);
    action
      matchtable_write_tunnel_lookup_miss(key, data);
    endaction
  endfunction

endinstance
interface TunnelLookupMiss;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkTunnelLookupMiss  (TunnelLookupMiss);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(31, 256, SizeOf#(TunnelLookupMissReqT), SizeOf#(TunnelLookupMissRspT)) matchTable <- mkMatchTable("tunnel_lookup_miss.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let i$p$v$6 = fromMaybe(?, meta.i$p$v$6);
    TunnelLookupMissReqT req = TunnelLookupMissReqT {i$p$v$4: i$p$v$4,i$p$v$6: i$p$v$6};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelLookupMissRspT resp = unpack(data);
      case (resp._action) matches
        NON_IP_TUNNEL_LOOKUP_MISS: begin
          BBRequest req = tagged NonIpTunnelLookupMissReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_TUNNEL_LOOKUP_MISS: begin
          BBRequest req = tagged Ipv4TunnelLookupMissReqT {pkt: pkt, l3_metadata$lkp_outer_l4_dport: l3_metadata$lkp_outer_l4_dport, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, ipv4$srcAddr: ipv4$srcAddr, ipv4$dstAddr: ipv4$dstAddr, ipv4$ttl: ipv4$ttl, ipv4$protocol: ipv4$protocol, l3_metadata$lkp_outer_l4_sport: l3_metadata$lkp_outer_l4_sport};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_TUNNEL_LOOKUP_MISS: begin
          BBRequest req = tagged Ipv6TunnelLookupMissReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, ipv6$srcAddr: ipv6$srcAddr, l3_metadata$lkp_outer_l4_dport: l3_metadata$lkp_outer_l4_dport, ipv6$dstAddr: ipv6$dstAddr, ipv6$hopLimit: ipv6$hopLimit, ipv6$nextHdr: ipv6$nextHdr, l3_metadata$lkp_outer_l4_sport: l3_metadata$lkp_outer_l4_sport};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NonIpTunnelLookupMissRspT {pkt: .pkt, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged TunnelLookupMissNonIpTunnelLookupMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4TunnelLookupMissRspT {pkt: .pkt, l3_metadata$lkp_ip_ttl: .l3_metadata$lkp_ip_ttl, ipv4_metadata$lkp_ipv4_da: .ipv4_metadata$lkp_ipv4_da, ipv4_metadata$lkp_ipv4_sa: .ipv4_metadata$lkp_ipv4_sa, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l3_metadata$lkp_l4_dport: .l3_metadata$lkp_l4_dport, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_sport: .l3_metadata$lkp_l4_sport, l3_metadata$lkp_ip_proto: .l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l3_metadata$lkp_ip_ttl = tagged Valid l3_metadata$lkp_ip_ttl;
        meta.ipv4_metadata$lkp_ipv4_da = tagged Valid ipv4_metadata$lkp_ipv4_da;
        meta.ipv4_metadata$lkp_ipv4_sa = tagged Valid ipv4_metadata$lkp_ipv4_sa;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l3_metadata$lkp_l4_dport = tagged Valid l3_metadata$lkp_l4_dport;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$lkp_l4_sport = tagged Valid l3_metadata$lkp_l4_sport;
        meta.l3_metadata$lkp_ip_proto = tagged Valid l3_metadata$lkp_ip_proto;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged TunnelLookupMissIpv4TunnelLookupMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6TunnelLookupMissRspT {pkt: .pkt, ipv6_metadata$lkp_ipv6_sa: .ipv6_metadata$lkp_ipv6_sa, ipv6_metadata$lkp_ipv6_da: .ipv6_metadata$lkp_ipv6_da, l3_metadata$lkp_l4_sport: .l3_metadata$lkp_l4_sport, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l3_metadata$lkp_ip_ttl: .l3_metadata$lkp_ip_ttl, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_dport: .l3_metadata$lkp_l4_dport, l3_metadata$lkp_ip_proto: .l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.ipv6_metadata$lkp_ipv6_sa = tagged Valid ipv6_metadata$lkp_ipv6_sa;
        meta.ipv6_metadata$lkp_ipv6_da = tagged Valid ipv6_metadata$lkp_ipv6_da;
        meta.l3_metadata$lkp_l4_sport = tagged Valid l3_metadata$lkp_l4_sport;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l3_metadata$lkp_ip_ttl = tagged Valid l3_metadata$lkp_ip_ttl;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$lkp_l4_dport = tagged Valid l3_metadata$lkp_l4_dport;
        meta.l3_metadata$lkp_ip_proto = tagged Valid l3_metadata$lkp_ip_proto;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged TunnelLookupMissIpv6TunnelLookupMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== TUNNEL_MISS ======

typedef struct {
  Bit#(7) padding;
  Bit#(Bool) valid_ipv4;
  Bit#(Bool) valid_ipv6;
} TunnelMissReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_MISS,
  NON_IP_TUNNEL_LOOKUP_MISS,
  IPV4_TUNNEL_LOOKUP_MISS,
  IPV6_TUNNEL_LOOKUP_MISS
} TunnelMissActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelMissActionT _action;
} TunnelMissRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_tunnel_miss(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_tunnel_miss(Bit#(9) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(30, 9, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(30) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_tunnel_miss(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(30) id, Bit#(9) key, Bit#(2) data);
    action
      matchtable_write_tunnel_miss(key, data);
    endaction
  endfunction

endinstance
interface TunnelMiss;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkTunnelMiss  (TunnelMiss);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(30, 256, SizeOf#(TunnelMissReqT), SizeOf#(TunnelMissRspT)) matchTable <- mkMatchTable("tunnel_miss.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let i$p$v$6 = fromMaybe(?, meta.i$p$v$6);
    TunnelMissReqT req = TunnelMissReqT {i$p$v$4: i$p$v$4,i$p$v$6: i$p$v$6};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelMissRspT resp = unpack(data);
      case (resp._action) matches
        NON_IP_TUNNEL_LOOKUP_MISS: begin
          BBRequest req = tagged NonIpTunnelLookupMissReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_TUNNEL_LOOKUP_MISS: begin
          BBRequest req = tagged Ipv4TunnelLookupMissReqT {pkt: pkt, l3_metadata$lkp_outer_l4_dport: l3_metadata$lkp_outer_l4_dport, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, ipv4$srcAddr: ipv4$srcAddr, ipv4$dstAddr: ipv4$dstAddr, ipv4$ttl: ipv4$ttl, ipv4$protocol: ipv4$protocol, l3_metadata$lkp_outer_l4_sport: l3_metadata$lkp_outer_l4_sport};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_TUNNEL_LOOKUP_MISS: begin
          BBRequest req = tagged Ipv6TunnelLookupMissReqT {pkt: pkt, ethernet$srcAddr: ethernet$srcAddr, ethernet$dstAddr: ethernet$dstAddr, ipv6$srcAddr: ipv6$srcAddr, l3_metadata$lkp_outer_l4_dport: l3_metadata$lkp_outer_l4_dport, ipv6$dstAddr: ipv6$dstAddr, ipv6$hopLimit: ipv6$hopLimit, ipv6$nextHdr: ipv6$nextHdr, l3_metadata$lkp_outer_l4_sport: l3_metadata$lkp_outer_l4_sport};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NonIpTunnelLookupMissRspT {pkt: .pkt, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged TunnelMissNonIpTunnelLookupMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4TunnelLookupMissRspT {pkt: .pkt, l3_metadata$lkp_ip_ttl: .l3_metadata$lkp_ip_ttl, ipv4_metadata$lkp_ipv4_da: .ipv4_metadata$lkp_ipv4_da, ipv4_metadata$lkp_ipv4_sa: .ipv4_metadata$lkp_ipv4_sa, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l3_metadata$lkp_l4_dport: .l3_metadata$lkp_l4_dport, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_sport: .l3_metadata$lkp_l4_sport, l3_metadata$lkp_ip_proto: .l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.l3_metadata$lkp_ip_ttl = tagged Valid l3_metadata$lkp_ip_ttl;
        meta.ipv4_metadata$lkp_ipv4_da = tagged Valid ipv4_metadata$lkp_ipv4_da;
        meta.ipv4_metadata$lkp_ipv4_sa = tagged Valid ipv4_metadata$lkp_ipv4_sa;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l3_metadata$lkp_l4_dport = tagged Valid l3_metadata$lkp_l4_dport;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$lkp_l4_sport = tagged Valid l3_metadata$lkp_l4_sport;
        meta.l3_metadata$lkp_ip_proto = tagged Valid l3_metadata$lkp_ip_proto;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged TunnelMissIpv4TunnelLookupMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6TunnelLookupMissRspT {pkt: .pkt, ipv6_metadata$lkp_ipv6_sa: .ipv6_metadata$lkp_ipv6_sa, ipv6_metadata$lkp_ipv6_da: .ipv6_metadata$lkp_ipv6_da, l3_metadata$lkp_l4_sport: .l3_metadata$lkp_l4_sport, intrinsic_metadata$mcast_grp: .intrinsic_metadata$mcast_grp, l3_metadata$lkp_ip_ttl: .l3_metadata$lkp_ip_ttl, l2_metadata$lkp_mac_sa: .l2_metadata$lkp_mac_sa, l3_metadata$lkp_l4_dport: .l3_metadata$lkp_l4_dport, l3_metadata$lkp_ip_proto: .l3_metadata$lkp_ip_proto, l2_metadata$lkp_mac_da: .l2_metadata$lkp_mac_da}: begin
        meta.ipv6_metadata$lkp_ipv6_sa = tagged Valid ipv6_metadata$lkp_ipv6_sa;
        meta.ipv6_metadata$lkp_ipv6_da = tagged Valid ipv6_metadata$lkp_ipv6_da;
        meta.l3_metadata$lkp_l4_sport = tagged Valid l3_metadata$lkp_l4_sport;
        meta.intrinsic_metadata$mcast_grp = tagged Valid intrinsic_metadata$mcast_grp;
        meta.l3_metadata$lkp_ip_ttl = tagged Valid l3_metadata$lkp_ip_ttl;
        meta.l2_metadata$lkp_mac_sa = tagged Valid l2_metadata$lkp_mac_sa;
        meta.l3_metadata$lkp_l4_dport = tagged Valid l3_metadata$lkp_l4_dport;
        meta.l3_metadata$lkp_ip_proto = tagged Valid l3_metadata$lkp_ip_proto;
        meta.l2_metadata$lkp_mac_da = tagged Valid l2_metadata$lkp_mac_da;
        MetadataResponse rsp = tagged TunnelMissIpv6TunnelLookupMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== URPF_BD ======

typedef struct {
  Bit#(4) padding;
  Bit#(16) l3_metadata$urpf_bd_group;
  Bit#(16) ingress_metadata$bd;
} UrpfBdReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_URPF_BD,
  NOP,
  URPF_BD_MISS
} UrpfBdActionT deriving (Bits, Eq, FShow);
typedef struct {
  UrpfBdActionT _action;
} UrpfBdRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_urpf_bd(Bit#(36) msgtype);
import "BDPI" function Action matchtable_write_urpf_bd(Bit#(36) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(13, 36, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(13) id, Bit#(36) key);
    actionvalue
      let v <- matchtable_read_urpf_bd(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(13) id, Bit#(36) key, Bit#(2) data);
    action
      matchtable_write_urpf_bd(key, data);
    endaction
  endfunction

endinstance
interface UrpfBd;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkUrpfBd  (UrpfBd);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(13, 1024, SizeOf#(UrpfBdReqT), SizeOf#(UrpfBdRspT)) matchTable <- mkMatchTable("urpf_bd.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$urpf_bd_group = fromMaybe(?, meta.l3_metadata$urpf_bd_group);
    let ingress_metadata$bd = fromMaybe(?, meta.ingress_metadata$bd);
    UrpfBdReqT req = UrpfBdReqT {l3_metadata$urpf_bd_group: l3_metadata$urpf_bd_group,ingress_metadata$bd: ingress_metadata$bd};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      UrpfBdRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        URPF_BD_MISS: begin
          BBRequest req = tagged UrpfBdMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged UrpfBdNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged UrpfBdMissRspT {pkt: .pkt, l3_metadata$urpf_check_fail: .l3_metadata$urpf_check_fail}: begin
        meta.l3_metadata$urpf_check_fail = tagged Valid l3_metadata$urpf_check_fail;
        MetadataResponse rsp = tagged UrpfBdUrpfBdMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== VALIDATE_MPLS_PACKET ======

typedef struct {
  Bit#(6) padding;
  Bit#(20) mpls0$label;
  Bit#(1) mpls0$bos;
  Bit#(Bool) valid_mpls0;
  Bit#(20) mpls1$label;
  Bit#(1) mpls1$bos;
  Bit#(Bool) valid_mpls1;
  Bit#(20) mpls2$label;
  Bit#(1) mpls2$bos;
  Bit#(Bool) valid_mpls2;
} ValidateMplsPacketReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_VALIDATE_MPLS_PACKET,
  SET_VALID_MPLS_LABEL1,
  SET_VALID_MPLS_LABEL2,
  SET_VALID_MPLS_LABEL3
} ValidateMplsPacketActionT deriving (Bits, Eq, FShow);
typedef struct {
  ValidateMplsPacketActionT _action;
} ValidateMplsPacketRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_validate_mpls_packet(Bit#(72) msgtype);
import "BDPI" function Action matchtable_write_validate_mpls_packet(Bit#(72) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(32, 72, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(32) id, Bit#(72) key);
    actionvalue
      let v <- matchtable_read_validate_mpls_packet(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(32) id, Bit#(72) key, Bit#(2) data);
    action
      matchtable_write_validate_mpls_packet(key, data);
    endaction
  endfunction

endinstance
interface ValidateMplsPacket;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkValidateMplsPacket  (ValidateMplsPacket);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(32, 512, SizeOf#(ValidateMplsPacketReqT), SizeOf#(ValidateMplsPacketRspT)) matchTable <- mkMatchTable("validate_mpls_packet.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let mpls0$label = fromMaybe(?, meta.mpls0$label);
    let mpls0$bos = fromMaybe(?, meta.mpls0$bos);
    let m$p$l$s$$0$ = fromMaybe(?, meta.m$p$l$s$$0$);
    let mpls1$label = fromMaybe(?, meta.mpls1$label);
    let mpls1$bos = fromMaybe(?, meta.mpls1$bos);
    let m$p$l$s$$1$ = fromMaybe(?, meta.m$p$l$s$$1$);
    let mpls2$label = fromMaybe(?, meta.mpls2$label);
    let mpls2$bos = fromMaybe(?, meta.mpls2$bos);
    let m$p$l$s$$2$ = fromMaybe(?, meta.m$p$l$s$$2$);
    ValidateMplsPacketReqT req = ValidateMplsPacketReqT {mpls0$label: mpls0$label,mpls0$bos: mpls0$bos,m$p$l$s$$0$: m$p$l$s$$0$,mpls1$label: mpls1$label,mpls1$bos: mpls1$bos,m$p$l$s$$1$: m$p$l$s$$1$,mpls2$label: mpls2$label,mpls2$bos: mpls2$bos,m$p$l$s$$2$: m$p$l$s$$2$};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ValidateMplsPacketRspT resp = unpack(data);
      case (resp._action) matches
        SET_VALID_MPLS_LABEL1: begin
          BBRequest req = tagged SetValidMplsLabel1ReqT {pkt: pkt, mpls0$exp: mpls0$exp, mpls0$label: mpls0$label};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_MPLS_LABEL2: begin
          BBRequest req = tagged SetValidMplsLabel2ReqT {pkt: pkt, mpls1$label: mpls1$label, mpls1$exp: mpls1$exp};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_MPLS_LABEL3: begin
          BBRequest req = tagged SetValidMplsLabel3ReqT {pkt: pkt, mpls2$label: mpls2$label, mpls2$exp: mpls2$exp};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetValidMplsLabel1RspT {pkt: .pkt, tunnel_metadata$mpls_label: .tunnel_metadata$mpls_label, tunnel_metadata$mpls_exp: .tunnel_metadata$mpls_exp}: begin
        meta.tunnel_metadata$mpls_label = tagged Valid tunnel_metadata$mpls_label;
        meta.tunnel_metadata$mpls_exp = tagged Valid tunnel_metadata$mpls_exp;
        MetadataResponse rsp = tagged ValidateMplsPacketSetValidMplsLabel1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidMplsLabel2RspT {pkt: .pkt, tunnel_metadata$mpls_label: .tunnel_metadata$mpls_label, tunnel_metadata$mpls_exp: .tunnel_metadata$mpls_exp}: begin
        meta.tunnel_metadata$mpls_label = tagged Valid tunnel_metadata$mpls_label;
        meta.tunnel_metadata$mpls_exp = tagged Valid tunnel_metadata$mpls_exp;
        MetadataResponse rsp = tagged ValidateMplsPacketSetValidMplsLabel2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidMplsLabel3RspT {pkt: .pkt, tunnel_metadata$mpls_label: .tunnel_metadata$mpls_label, tunnel_metadata$mpls_exp: .tunnel_metadata$mpls_exp}: begin
        meta.tunnel_metadata$mpls_label = tagged Valid tunnel_metadata$mpls_label;
        meta.tunnel_metadata$mpls_exp = tagged Valid tunnel_metadata$mpls_exp;
        MetadataResponse rsp = tagged ValidateMplsPacketSetValidMplsLabel3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== VALIDATE_OUTER_ETHERNET ======

typedef struct {
  Bit#(1) padding;
  Bit#(48) ethernet$srcAddr;
  Bit#(48) ethernet$dstAddr;
  Bit#(Bool) valid_vlan_tag_0;
  Bit#(Bool) valid_vlan_tag_1;
} ValidateOuterEthernetReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_VALIDATE_OUTER_ETHERNET,
  MALFORMED_OUTER_ETHERNET_PACKET,
  SET_VALID_OUTER_UNICAST_PACKET_UNTAGGED,
  SET_VALID_OUTER_UNICAST_PACKET_SINGLE_TAGGED,
  SET_VALID_OUTER_UNICAST_PACKET_DOUBLE_TAGGED,
  SET_VALID_OUTER_UNICAST_PACKET_QINQ_TAGGED,
  SET_VALID_OUTER_MULTICAST_PACKET_UNTAGGED,
  SET_VALID_OUTER_MULTICAST_PACKET_SINGLE_TAGGED,
  SET_VALID_OUTER_MULTICAST_PACKET_DOUBLE_TAGGED,
  SET_VALID_OUTER_MULTICAST_PACKET_QINQ_TAGGED,
  SET_VALID_OUTER_BROADCAST_PACKET_UNTAGGED,
  SET_VALID_OUTER_BROADCAST_PACKET_SINGLE_TAGGED,
  SET_VALID_OUTER_BROADCAST_PACKET_DOUBLE_TAGGED,
  SET_VALID_OUTER_BROADCAST_PACKET_QINQ_TAGGED
} ValidateOuterEthernetActionT deriving (Bits, Eq, FShow);
typedef struct {
  ValidateOuterEthernetActionT _action;
  Bit#(8) runtime_drop_reason;
} ValidateOuterEthernetRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(12)) matchtable_read_validate_outer_ethernet(Bit#(99) msgtype);
import "BDPI" function Action matchtable_write_validate_outer_ethernet(Bit#(99) msgtype, Bit#(12) data);
`endif
instance MatchTableSim#(1, 99, 12);
  function ActionValue#(Bit#(12)) matchtable_read(Bit#(1) id, Bit#(99) key);
    actionvalue
      let v <- matchtable_read_validate_outer_ethernet(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(1) id, Bit#(99) key, Bit#(12) data);
    action
      matchtable_write_validate_outer_ethernet(key, data);
    endaction
  endfunction

endinstance
interface ValidateOuterEthernet;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
  interface Client #(BBRequest, BBResponse) next_control_state_9;
  interface Client #(BBRequest, BBResponse) next_control_state_10;
  interface Client #(BBRequest, BBResponse) next_control_state_11;
  interface Client #(BBRequest, BBResponse) next_control_state_12;
endinterface
(* synthesize *)
module mkValidateOuterEthernet  (ValidateOuterEthernet);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(13, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(13, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(1, 512, SizeOf#(ValidateOuterEthernetReqT), SizeOf#(ValidateOuterEthernetRspT)) matchTable <- mkMatchTable("validate_outer_ethernet.dat");
  Vector#(13, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(13) readyChannel = -1;
  for (Integer i=12; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ethernet$srcAddr = fromMaybe(?, meta.ethernet$srcAddr);
    let ethernet$dstAddr = fromMaybe(?, meta.ethernet$dstAddr);
    let v$l$a$n$_$t$a$g$_$$0$ = fromMaybe(?, meta.v$l$a$n$_$t$a$g$_$$0$);
    let v$l$a$n$_$t$a$g$_$$1$ = fromMaybe(?, meta.v$l$a$n$_$t$a$g$_$$1$);
    ValidateOuterEthernetReqT req = ValidateOuterEthernetReqT {ethernet$srcAddr: ethernet$srcAddr,ethernet$dstAddr: ethernet$dstAddr,v$l$a$n$_$t$a$g$_$$0$: v$l$a$n$_$t$a$g$_$$0$,v$l$a$n$_$t$a$g$_$$1$: v$l$a$n$_$t$a$g$_$$1$};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ValidateOuterEthernetRspT resp = unpack(data);
      case (resp._action) matches
        MALFORMED_OUTER_ETHERNET_PACKET: begin
          BBRequest req = tagged MalformedOuterEthernetPacketReqT {pkt: pkt, runtime_drop_reason: resp.runtime_drop_reason};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_UNICAST_PACKET_UNTAGGED: begin
          BBRequest req = tagged SetValidOuterUnicastPacketUntaggedReqT {pkt: pkt, ethernet$etherType: ethernet$etherType};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_UNICAST_PACKET_SINGLE_TAGGED: begin
          BBRequest req = tagged SetValidOuterUnicastPacketSingleTaggedReqT {pkt: pkt, vlan_tag_0$etherType: vlan_tag_0$etherType};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_UNICAST_PACKET_DOUBLE_TAGGED: begin
          BBRequest req = tagged SetValidOuterUnicastPacketDoubleTaggedReqT {pkt: pkt, vlan_tag_1$etherType: vlan_tag_1$etherType};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_UNICAST_PACKET_QINQ_TAGGED: begin
          BBRequest req = tagged SetValidOuterUnicastPacketQinqTaggedReqT {pkt: pkt, ethernet$etherType: ethernet$etherType};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_MULTICAST_PACKET_UNTAGGED: begin
          BBRequest req = tagged SetValidOuterMulticastPacketUntaggedReqT {pkt: pkt, ethernet$etherType: ethernet$etherType};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_MULTICAST_PACKET_SINGLE_TAGGED: begin
          BBRequest req = tagged SetValidOuterMulticastPacketSingleTaggedReqT {pkt: pkt, vlan_tag_0$etherType: vlan_tag_0$etherType};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_MULTICAST_PACKET_DOUBLE_TAGGED: begin
          BBRequest req = tagged SetValidOuterMulticastPacketDoubleTaggedReqT {pkt: pkt, vlan_tag_1$etherType: vlan_tag_1$etherType};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_MULTICAST_PACKET_QINQ_TAGGED: begin
          BBRequest req = tagged SetValidOuterMulticastPacketQinqTaggedReqT {pkt: pkt, ethernet$etherType: ethernet$etherType};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_BROADCAST_PACKET_UNTAGGED: begin
          BBRequest req = tagged SetValidOuterBroadcastPacketUntaggedReqT {pkt: pkt, ethernet$etherType: ethernet$etherType};
          bbReqFifo[9].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_BROADCAST_PACKET_SINGLE_TAGGED: begin
          BBRequest req = tagged SetValidOuterBroadcastPacketSingleTaggedReqT {pkt: pkt, vlan_tag_0$etherType: vlan_tag_0$etherType};
          bbReqFifo[10].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_BROADCAST_PACKET_DOUBLE_TAGGED: begin
          BBRequest req = tagged SetValidOuterBroadcastPacketDoubleTaggedReqT {pkt: pkt, vlan_tag_1$etherType: vlan_tag_1$etherType};
          bbReqFifo[11].enq(req); //FIXME: replace with RXTX.
        end
        SET_VALID_OUTER_BROADCAST_PACKET_QINQ_TAGGED: begin
          BBRequest req = tagged SetValidOuterBroadcastPacketQinqTaggedReqT {pkt: pkt, ethernet$etherType: ethernet$etherType};
          bbReqFifo[12].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged MalformedOuterEthernetPacketRspT {pkt: .pkt, ingress_metadata$drop_reason: .ingress_metadata$drop_reason, ingress_metadata$drop_flag: .ingress_metadata$drop_flag}: begin
        meta.ingress_metadata$drop_reason = tagged Valid ingress_metadata$drop_reason;
        meta.ingress_metadata$drop_flag = tagged Valid ingress_metadata$drop_flag;
        MetadataResponse rsp = tagged ValidateOuterEthernetMalformedOuterEthernetPacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterUnicastPacketUntaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterUnicastPacketUntaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterUnicastPacketSingleTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterUnicastPacketSingleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterUnicastPacketDoubleTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterUnicastPacketDoubleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterUnicastPacketQinqTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterUnicastPacketQinqTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterMulticastPacketUntaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterMulticastPacketUntaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterMulticastPacketSingleTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterMulticastPacketSingleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterMulticastPacketDoubleTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterMulticastPacketDoubleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterMulticastPacketQinqTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterMulticastPacketQinqTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterBroadcastPacketUntaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterBroadcastPacketUntaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterBroadcastPacketSingleTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterBroadcastPacketSingleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterBroadcastPacketDoubleTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterBroadcastPacketDoubleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetValidOuterBroadcastPacketQinqTaggedRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$lkp_mac_type: .l2_metadata$lkp_mac_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$lkp_mac_type = tagged Valid l2_metadata$lkp_mac_type;
        MetadataResponse rsp = tagged ValidateOuterEthernetSetValidOuterBroadcastPacketQinqTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
  interface next_control_state_9 = toClient(bbReqFifo[9], bbRspFifo[9]);
  interface next_control_state_10 = toClient(bbReqFifo[10], bbRspFifo[10]);
  interface next_control_state_11 = toClient(bbReqFifo[11], bbRspFifo[11]);
  interface next_control_state_12 = toClient(bbReqFifo[12], bbRspFifo[12]);
endmodule

// ====== VALIDATE_OUTER_IPV4_PACKET ======

typedef struct {
  Bit#(1) padding;
  Bit#(4) ipv4$version;
  Bit#(8) ipv4$ttl;
  Bit#(32) ipv4$srcAddr;
} ValidateOuterIpv4PacketReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_VALIDATE_OUTER_IPV4_PACKET,
  SET_VALID_OUTER_IPV4_PACKET,
  SET_MALFORMED_OUTER_IPV4_PACKET
} ValidateOuterIpv4PacketActionT deriving (Bits, Eq, FShow);
typedef struct {
  ValidateOuterIpv4PacketActionT _action;
  Bit#(8) runtime_drop_reason;
} ValidateOuterIpv4PacketRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(10)) matchtable_read_validate_outer_ipv4_packet(Bit#(45) msgtype);
import "BDPI" function Action matchtable_write_validate_outer_ipv4_packet(Bit#(45) msgtype, Bit#(10) data);
`endif
instance MatchTableSim#(14, 45, 10);
  function ActionValue#(Bit#(10)) matchtable_read(Bit#(14) id, Bit#(45) key);
    actionvalue
      let v <- matchtable_read_validate_outer_ipv4_packet(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(14) id, Bit#(45) key, Bit#(10) data);
    action
      matchtable_write_validate_outer_ipv4_packet(key, data);
    endaction
  endfunction

endinstance
interface ValidateOuterIpv4Packet;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkValidateOuterIpv4Packet  (ValidateOuterIpv4Packet);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(14, 512, SizeOf#(ValidateOuterIpv4PacketReqT), SizeOf#(ValidateOuterIpv4PacketRspT)) matchTable <- mkMatchTable("validate_outer_ipv4_packet.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ipv4$version = fromMaybe(?, meta.ipv4$version);
    let ipv4$ttl = fromMaybe(?, meta.ipv4$ttl);
    let ipv4$srcAddr = fromMaybe(?, meta.ipv4$srcAddr);
    ValidateOuterIpv4PacketReqT req = ValidateOuterIpv4PacketReqT {ipv4$version: ipv4$version,ipv4$ttl: ipv4$ttl,ipv4$srcAddr: ipv4$srcAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ValidateOuterIpv4PacketRspT resp = unpack(data);
      case (resp._action) matches
        SET_VALID_OUTER_IPV4_PACKET: begin
          BBRequest req = tagged SetValidOuterIpv4PacketReqT {pkt: pkt, ipv4$diffserv: ipv4$diffserv, ipv4$version: ipv4$version};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_MALFORMED_OUTER_IPV4_PACKET: begin
          BBRequest req = tagged SetMalformedOuterIpv4PacketReqT {pkt: pkt, runtime_drop_reason: resp.runtime_drop_reason};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetValidOuterIpv4PacketRspT {pkt: .pkt, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, l3_metadata$lkp_ip_version: .l3_metadata$lkp_ip_version}: begin
        meta.l3_metadata$lkp_ip_tc = tagged Valid l3_metadata$lkp_ip_tc;
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.l3_metadata$lkp_ip_version = tagged Valid l3_metadata$lkp_ip_version;
        MetadataResponse rsp = tagged ValidateOuterIpv4PacketSetValidOuterIpv4PacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMalformedOuterIpv4PacketRspT {pkt: .pkt, ingress_metadata$drop_reason: .ingress_metadata$drop_reason, ingress_metadata$drop_flag: .ingress_metadata$drop_flag}: begin
        meta.ingress_metadata$drop_reason = tagged Valid ingress_metadata$drop_reason;
        meta.ingress_metadata$drop_flag = tagged Valid ingress_metadata$drop_flag;
        MetadataResponse rsp = tagged ValidateOuterIpv4PacketSetMalformedOuterIpv4PacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== VALIDATE_OUTER_IPV6_PACKET ======

typedef struct {
  Bit#(4) padding;
  Bit#(4) ipv6$version;
  Bit#(8) ipv6$hopLimit;
  Bit#(128) ipv6$srcAddr;
} ValidateOuterIpv6PacketReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_VALIDATE_OUTER_IPV6_PACKET,
  SET_VALID_OUTER_IPV6_PACKET,
  SET_MALFORMED_OUTER_IPV6_PACKET
} ValidateOuterIpv6PacketActionT deriving (Bits, Eq, FShow);
typedef struct {
  ValidateOuterIpv6PacketActionT _action;
  Bit#(8) runtime_drop_reason;
} ValidateOuterIpv6PacketRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(10)) matchtable_read_validate_outer_ipv6_packet(Bit#(144) msgtype);
import "BDPI" function Action matchtable_write_validate_outer_ipv6_packet(Bit#(144) msgtype, Bit#(10) data);
`endif
instance MatchTableSim#(19, 144, 10);
  function ActionValue#(Bit#(10)) matchtable_read(Bit#(19) id, Bit#(144) key);
    actionvalue
      let v <- matchtable_read_validate_outer_ipv6_packet(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(19) id, Bit#(144) key, Bit#(10) data);
    action
      matchtable_write_validate_outer_ipv6_packet(key, data);
    endaction
  endfunction

endinstance
interface ValidateOuterIpv6Packet;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkValidateOuterIpv6Packet  (ValidateOuterIpv6Packet);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(19, 512, SizeOf#(ValidateOuterIpv6PacketReqT), SizeOf#(ValidateOuterIpv6PacketRspT)) matchTable <- mkMatchTable("validate_outer_ipv6_packet.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let ipv6$version = fromMaybe(?, meta.ipv6$version);
    let ipv6$hopLimit = fromMaybe(?, meta.ipv6$hopLimit);
    let ipv6$srcAddr = fromMaybe(?, meta.ipv6$srcAddr);
    ValidateOuterIpv6PacketReqT req = ValidateOuterIpv6PacketReqT {ipv6$version: ipv6$version,ipv6$hopLimit: ipv6$hopLimit,ipv6$srcAddr: ipv6$srcAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ValidateOuterIpv6PacketRspT resp = unpack(data);
      case (resp._action) matches
        SET_VALID_OUTER_IPV6_PACKET: begin
          BBRequest req = tagged SetValidOuterIpv6PacketReqT {pkt: pkt, ipv6$version: ipv6$version, ipv6$trafficClass: ipv6$trafficClass};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_MALFORMED_OUTER_IPV6_PACKET: begin
          BBRequest req = tagged SetMalformedOuterIpv6PacketReqT {pkt: pkt, runtime_drop_reason: resp.runtime_drop_reason};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetValidOuterIpv6PacketRspT {pkt: .pkt, l3_metadata$lkp_ip_tc: .l3_metadata$lkp_ip_tc, l3_metadata$lkp_ip_type: .l3_metadata$lkp_ip_type, l3_metadata$lkp_ip_version: .l3_metadata$lkp_ip_version}: begin
        meta.l3_metadata$lkp_ip_tc = tagged Valid l3_metadata$lkp_ip_tc;
        meta.l3_metadata$lkp_ip_type = tagged Valid l3_metadata$lkp_ip_type;
        meta.l3_metadata$lkp_ip_version = tagged Valid l3_metadata$lkp_ip_version;
        MetadataResponse rsp = tagged ValidateOuterIpv6PacketSetValidOuterIpv6PacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMalformedOuterIpv6PacketRspT {pkt: .pkt, ingress_metadata$drop_reason: .ingress_metadata$drop_reason, ingress_metadata$drop_flag: .ingress_metadata$drop_flag}: begin
        meta.ingress_metadata$drop_reason = tagged Valid ingress_metadata$drop_reason;
        meta.ingress_metadata$drop_flag = tagged Valid ingress_metadata$drop_flag;
        MetadataResponse rsp = tagged ValidateOuterIpv6PacketSetMalformedOuterIpv6PacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== VALIDATE_PACKET ======

typedef struct {
  Bit#(48) l2_metadata$lkp_mac_sa;
  Bit#(48) l2_metadata$lkp_mac_da;
  Bit#(2) l3_metadata$lkp_ip_type;
  Bit#(8) l3_metadata$lkp_ip_ttl;
  Bit#(4) l3_metadata$lkp_ip_version;
  Bit#(32) ipv4_metadata$lkp_ipv4_sa;
  Bit#(128) ipv6_metadata$lkp_ipv6_sa;
} ValidatePacketReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_VALIDATE_PACKET,
  NOP,
  SET_UNICAST,
  SET_UNICAST_AND_IPV6_SRC_IS_LINK_LOCAL,
  SET_MULTICAST,
  SET_MULTICAST_AND_IPV6_SRC_IS_LINK_LOCAL,
  SET_BROADCAST,
  SET_MALFORMED_PACKET
} ValidatePacketActionT deriving (Bits, Eq, FShow);
typedef struct {
  ValidatePacketActionT _action;
  Bit#(8) runtime_drop_reason;
} ValidatePacketRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(11)) matchtable_read_validate_packet(Bit#(270) msgtype);
import "BDPI" function Action matchtable_write_validate_packet(Bit#(270) msgtype, Bit#(11) data);
`endif
instance MatchTableSim#(11, 270, 11);
  function ActionValue#(Bit#(11)) matchtable_read(Bit#(11) id, Bit#(270) key);
    actionvalue
      let v <- matchtable_read_validate_packet(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(11) id, Bit#(270) key, Bit#(11) data);
    action
      matchtable_write_validate_packet(key, data);
    endaction
  endfunction

endinstance
interface ValidatePacket;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
endinterface
(* synthesize *)
module mkValidatePacket  (ValidatePacket);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(7, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(7, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(11, 512, SizeOf#(ValidatePacketReqT), SizeOf#(ValidatePacketRspT)) matchTable <- mkMatchTable("validate_packet.dat");
  Vector#(7, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(7) readyChannel = -1;
  for (Integer i=6; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l2_metadata$lkp_mac_sa = fromMaybe(?, meta.l2_metadata$lkp_mac_sa);
    let l2_metadata$lkp_mac_da = fromMaybe(?, meta.l2_metadata$lkp_mac_da);
    let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
    let l3_metadata$lkp_ip_ttl = fromMaybe(?, meta.l3_metadata$lkp_ip_ttl);
    let l3_metadata$lkp_ip_version = fromMaybe(?, meta.l3_metadata$lkp_ip_version);
    let ipv4_metadata$lkp_ipv4_sa = fromMaybe(?, meta.ipv4_metadata$lkp_ipv4_sa);
    let ipv6_metadata$lkp_ipv6_sa = fromMaybe(?, meta.ipv6_metadata$lkp_ipv6_sa);
    ValidatePacketReqT req = ValidatePacketReqT {l2_metadata$lkp_mac_sa: l2_metadata$lkp_mac_sa,l2_metadata$lkp_mac_da: l2_metadata$lkp_mac_da,l3_metadata$lkp_ip_type: l3_metadata$lkp_ip_type,l3_metadata$lkp_ip_ttl: l3_metadata$lkp_ip_ttl,l3_metadata$lkp_ip_version: l3_metadata$lkp_ip_version,ipv4_metadata$lkp_ipv4_sa: ipv4_metadata$lkp_ipv4_sa,ipv6_metadata$lkp_ipv6_sa: ipv6_metadata$lkp_ipv6_sa};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ValidatePacketRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_UNICAST: begin
          BBRequest req = tagged SetUnicastReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_UNICAST_AND_IPV6_SRC_IS_LINK_LOCAL: begin
          BBRequest req = tagged SetUnicastAndIpv6SrcIsLinkLocalReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        SET_MULTICAST: begin
          BBRequest req = tagged SetMulticastReqT {pkt: pkt};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        SET_MULTICAST_AND_IPV6_SRC_IS_LINK_LOCAL: begin
          BBRequest req = tagged SetMulticastAndIpv6SrcIsLinkLocalReqT {pkt: pkt};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        SET_BROADCAST: begin
          BBRequest req = tagged SetBroadcastReqT {pkt: pkt};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        SET_MALFORMED_PACKET: begin
          BBRequest req = tagged SetMalformedPacketReqT {pkt: pkt, runtime_drop_reason: resp.runtime_drop_reason};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged ValidatePacketNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetUnicastRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        MetadataResponse rsp = tagged ValidatePacketSetUnicastRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetUnicastAndIpv6SrcIsLinkLocalRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, ipv6_metadata$ipv6_src_is_link_local: .ipv6_metadata$ipv6_src_is_link_local}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.ipv6_metadata$ipv6_src_is_link_local = tagged Valid ipv6_metadata$ipv6_src_is_link_local;
        MetadataResponse rsp = tagged ValidatePacketSetUnicastAndIpv6SrcIsLinkLocalRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMulticastRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$bd_stats_idx: .l2_metadata$bd_stats_idx}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$bd_stats_idx = tagged Valid l2_metadata$bd_stats_idx;
        MetadataResponse rsp = tagged ValidatePacketSetMulticastRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMulticastAndIpv6SrcIsLinkLocalRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, ipv6_metadata$ipv6_src_is_link_local: .ipv6_metadata$ipv6_src_is_link_local, l2_metadata$bd_stats_idx: .l2_metadata$bd_stats_idx}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.ipv6_metadata$ipv6_src_is_link_local = tagged Valid ipv6_metadata$ipv6_src_is_link_local;
        meta.l2_metadata$bd_stats_idx = tagged Valid l2_metadata$bd_stats_idx;
        MetadataResponse rsp = tagged ValidatePacketSetMulticastAndIpv6SrcIsLinkLocalRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetBroadcastRspT {pkt: .pkt, l2_metadata$lkp_pkt_type: .l2_metadata$lkp_pkt_type, l2_metadata$bd_stats_idx: .l2_metadata$bd_stats_idx}: begin
        meta.l2_metadata$lkp_pkt_type = tagged Valid l2_metadata$lkp_pkt_type;
        meta.l2_metadata$bd_stats_idx = tagged Valid l2_metadata$bd_stats_idx;
        MetadataResponse rsp = tagged ValidatePacketSetBroadcastRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMalformedPacketRspT {pkt: .pkt, ingress_metadata$drop_reason: .ingress_metadata$drop_reason, ingress_metadata$drop_flag: .ingress_metadata$drop_flag}: begin
        meta.ingress_metadata$drop_reason = tagged Valid ingress_metadata$drop_reason;
        meta.ingress_metadata$drop_flag = tagged Valid ingress_metadata$drop_flag;
        MetadataResponse rsp = tagged ValidatePacketSetMalformedPacketRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
endmodule

// ====== INGRESS ======

interface Ingress;
  interface Client#(MetadataRequest, MetadataResponse) next;
endinterface
module mkIngress #(Vector#(numClients, Client#(MetadataRequest, MetadataResponse)) mdc) (Ingress);
  FIFOF#(MetadataRequest) default_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) default_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) acl_stats_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) acl_stats_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) bd_flood_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) bd_flood_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) compute_ipv4_hashes_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) compute_ipv4_hashes_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) compute_ipv6_hashes_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) compute_ipv6_hashes_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) compute_non_ip_hashes_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) compute_non_ip_hashes_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) compute_other_hashes_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) compute_other_hashes_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) dmac_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) dmac_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) drop_stats_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) drop_stats_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ecmp_group_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ecmp_group_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) fabric_ingress_dst_lkp_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) fabric_ingress_dst_lkp_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) fabric_ingress_src_lkp_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) fabric_ingress_src_lkp_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) fabric_lag_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) fabric_lag_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) fwd_result_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) fwd_result_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ingress_bd_stats_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ingress_bd_stats_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ingress_port_mapping_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ingress_port_mapping_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ingress_port_properties_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ingress_port_properties_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_sink_update_outer_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_sink_update_outer_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_source_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_source_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_terminate_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_terminate_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ip_acl_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ip_acl_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipsg_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipsg_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipsg_permit_special_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipsg_permit_special_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_dest_vtep_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_dest_vtep_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_fib_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_fib_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_fib_lpm_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_fib_lpm_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_multicast_bridge_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_multicast_bridge_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_multicast_bridge_star_g_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_multicast_bridge_star_g_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_multicast_route_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_multicast_route_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_multicast_route_star_g_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_multicast_route_star_g_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_racl_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_racl_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_src_vtep_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_src_vtep_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_urpf_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_urpf_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv4_urpf_lpm_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv4_urpf_lpm_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_acl_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_acl_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_dest_vtep_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_dest_vtep_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_fib_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_fib_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_fib_lpm_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_fib_lpm_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_multicast_bridge_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_multicast_bridge_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_multicast_bridge_star_g_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_multicast_bridge_star_g_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_multicast_route_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_multicast_route_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_multicast_route_star_g_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_multicast_route_star_g_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_racl_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_racl_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_src_vtep_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_src_vtep_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_urpf_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_urpf_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) ipv6_urpf_lpm_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) ipv6_urpf_lpm_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) lag_group_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) lag_group_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) learn_notify_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) learn_notify_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) mac_acl_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) mac_acl_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) meter_action_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) meter_action_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) meter_index_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) meter_index_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) mpls_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) mpls_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) native_packet_over_fabric_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) native_packet_over_fabric_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) nexthop_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) nexthop_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) outer_ipv4_multicast_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) outer_ipv4_multicast_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) outer_ipv4_multicast_star_g_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) outer_ipv4_multicast_star_g_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) outer_ipv6_multicast_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) outer_ipv6_multicast_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) outer_ipv6_multicast_star_g_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) outer_ipv6_multicast_star_g_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) outer_rmac_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) outer_rmac_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) port_vlan_mapping_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) port_vlan_mapping_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) qos_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) qos_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) rmac_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) rmac_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) sflow_ing_take_sample_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) sflow_ing_take_sample_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) sflow_ingress_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) sflow_ingress_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) smac_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) smac_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) spanning_tree_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) spanning_tree_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) storm_control_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) storm_control_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) storm_control_stats_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) storm_control_stats_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) switch_config_params_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) switch_config_params_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) system_acl_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) system_acl_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_lookup_miss_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_lookup_miss_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_miss_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_miss_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) urpf_bd_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) urpf_bd_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) validate_mpls_packet_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) validate_mpls_packet_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) validate_outer_ethernet_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) validate_outer_ethernet_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) validate_outer_ipv4_packet_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) validate_outer_ipv4_packet_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) validate_outer_ipv6_packet_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) validate_outer_ipv6_packet_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) validate_packet_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) validate_packet_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) next_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) next_rsp_ff <- mkFIFOF;
  Vector#(numClients, Server#(MetadataRequest, MetadataResponse)) mds = replicate(toServer(default_req_ff, default_rsp_ff));
  mkConnection(mds, mdc);
  AclStats acl_stats <- mkAclStats();
  BdFlood bd_flood <- mkBdFlood();
  ComputeIpv4Hashes compute_ipv4_hashes <- mkComputeIpv4Hashes();
  ComputeIpv6Hashes compute_ipv6_hashes <- mkComputeIpv6Hashes();
  ComputeNonIpHashes compute_non_ip_hashes <- mkComputeNonIpHashes();
  ComputeOtherHashes compute_other_hashes <- mkComputeOtherHashes();
  Dmac dmac <- mkDmac();
  DropStats drop_stats <- mkDropStats();
  EcmpGroup ecmp_group <- mkEcmpGroup();
  FabricIngressDstLkp fabric_ingress_dst_lkp <- mkFabricIngressDstLkp();
  FabricIngressSrcLkp fabric_ingress_src_lkp <- mkFabricIngressSrcLkp();
  FabricLag fabric_lag <- mkFabricLag();
  FwdResult fwd_result <- mkFwdResult();
  IngressBdStats ingress_bd_stats <- mkIngressBdStats();
  IngressPortMapping ingress_port_mapping <- mkIngressPortMapping();
  IngressPortProperties ingress_port_properties <- mkIngressPortProperties();
  IntSinkUpdateOuter int_sink_update_outer <- mkIntSinkUpdateOuter();
  IntSource int_source <- mkIntSource();
  IntTerminate int_terminate <- mkIntTerminate();
  IpAcl ip_acl <- mkIpAcl();
  Ipsg ipsg <- mkIpsg();
  IpsgPermitSpecial ipsg_permit_special <- mkIpsgPermitSpecial();
  Ipv4DestVtep ipv4_dest_vtep <- mkIpv4DestVtep();
  Ipv4Fib ipv4_fib <- mkIpv4Fib();
  Ipv4FibLpm ipv4_fib_lpm <- mkIpv4FibLpm();
  Ipv4MulticastBridge ipv4_multicast_bridge <- mkIpv4MulticastBridge();
  Ipv4MulticastBridgeStarG ipv4_multicast_bridge_star_g <- mkIpv4MulticastBridgeStarG();
  Ipv4MulticastRoute ipv4_multicast_route <- mkIpv4MulticastRoute();
  Ipv4MulticastRouteStarG ipv4_multicast_route_star_g <- mkIpv4MulticastRouteStarG();
  Ipv4Racl ipv4_racl <- mkIpv4Racl();
  Ipv4SrcVtep ipv4_src_vtep <- mkIpv4SrcVtep();
  Ipv4Urpf ipv4_urpf <- mkIpv4Urpf();
  Ipv4UrpfLpm ipv4_urpf_lpm <- mkIpv4UrpfLpm();
  Ipv6Acl ipv6_acl <- mkIpv6Acl();
  Ipv6DestVtep ipv6_dest_vtep <- mkIpv6DestVtep();
  Ipv6Fib ipv6_fib <- mkIpv6Fib();
  Ipv6FibLpm ipv6_fib_lpm <- mkIpv6FibLpm();
  Ipv6MulticastBridge ipv6_multicast_bridge <- mkIpv6MulticastBridge();
  Ipv6MulticastBridgeStarG ipv6_multicast_bridge_star_g <- mkIpv6MulticastBridgeStarG();
  Ipv6MulticastRoute ipv6_multicast_route <- mkIpv6MulticastRoute();
  Ipv6MulticastRouteStarG ipv6_multicast_route_star_g <- mkIpv6MulticastRouteStarG();
  Ipv6Racl ipv6_racl <- mkIpv6Racl();
  Ipv6SrcVtep ipv6_src_vtep <- mkIpv6SrcVtep();
  Ipv6Urpf ipv6_urpf <- mkIpv6Urpf();
  Ipv6UrpfLpm ipv6_urpf_lpm <- mkIpv6UrpfLpm();
  LagGroup lag_group <- mkLagGroup();
  LearnNotify learn_notify <- mkLearnNotify();
  MacAcl mac_acl <- mkMacAcl();
  MeterAction meter_action <- mkMeterAction();
  MeterIndex meter_index <- mkMeterIndex();
  Mpls mpls <- mkMpls();
  NativePacketOverFabric native_packet_over_fabric <- mkNativePacketOverFabric();
  Nexthop nexthop <- mkNexthop();
  OuterIpv4Multicast outer_ipv4_multicast <- mkOuterIpv4Multicast();
  OuterIpv4MulticastStarG outer_ipv4_multicast_star_g <- mkOuterIpv4MulticastStarG();
  OuterIpv6Multicast outer_ipv6_multicast <- mkOuterIpv6Multicast();
  OuterIpv6MulticastStarG outer_ipv6_multicast_star_g <- mkOuterIpv6MulticastStarG();
  OuterRmac outer_rmac <- mkOuterRmac();
  PortVlanMapping port_vlan_mapping <- mkPortVlanMapping();
  Qos qos <- mkQos();
  Rmac rmac <- mkRmac();
  SflowIngTakeSample sflow_ing_take_sample <- mkSflowIngTakeSample();
  SflowIngress sflow_ingress <- mkSflowIngress();
  Smac smac <- mkSmac();
  SpanningTree spanning_tree <- mkSpanningTree();
  StormControl storm_control <- mkStormControl();
  StormControlStats storm_control_stats <- mkStormControlStats();
  SwitchConfigParams switch_config_params <- mkSwitchConfigParams();
  SystemAcl system_acl <- mkSystemAcl();
  Tunnel tunnel <- mkTunnel();
  TunnelLookupMiss tunnel_lookup_miss <- mkTunnelLookupMiss();
  TunnelMiss tunnel_miss <- mkTunnelMiss();
  UrpfBd urpf_bd <- mkUrpfBd();
  ValidateMplsPacket validate_mpls_packet <- mkValidateMplsPacket();
  ValidateOuterEthernet validate_outer_ethernet <- mkValidateOuterEthernet();
  ValidateOuterIpv4Packet validate_outer_ipv4_packet <- mkValidateOuterIpv4Packet();
  ValidateOuterIpv6Packet validate_outer_ipv6_packet <- mkValidateOuterIpv6Packet();
  ValidatePacket validate_packet <- mkValidatePacket();
  mkConnection(toClient(acl_stats_req_ff, acl_stats_rsp_ff), acl_stats.prev_control_state_0);
  mkConnection(toClient(bd_flood_req_ff, bd_flood_rsp_ff), bd_flood.prev_control_state_0);
  mkConnection(toClient(compute_ipv4_hashes_req_ff, compute_ipv4_hashes_rsp_ff), compute_ipv4_hashes.prev_control_state_0);
  mkConnection(toClient(compute_ipv6_hashes_req_ff, compute_ipv6_hashes_rsp_ff), compute_ipv6_hashes.prev_control_state_0);
  mkConnection(toClient(compute_non_ip_hashes_req_ff, compute_non_ip_hashes_rsp_ff), compute_non_ip_hashes.prev_control_state_0);
  mkConnection(toClient(compute_other_hashes_req_ff, compute_other_hashes_rsp_ff), compute_other_hashes.prev_control_state_0);
  mkConnection(toClient(dmac_req_ff, dmac_rsp_ff), dmac.prev_control_state_0);
  mkConnection(toClient(drop_stats_req_ff, drop_stats_rsp_ff), drop_stats.prev_control_state_0);
  mkConnection(toClient(ecmp_group_req_ff, ecmp_group_rsp_ff), ecmp_group.prev_control_state_0);
  mkConnection(toClient(fabric_ingress_dst_lkp_req_ff, fabric_ingress_dst_lkp_rsp_ff), fabric_ingress_dst_lkp.prev_control_state_0);
  mkConnection(toClient(fabric_ingress_src_lkp_req_ff, fabric_ingress_src_lkp_rsp_ff), fabric_ingress_src_lkp.prev_control_state_0);
  mkConnection(toClient(fabric_lag_req_ff, fabric_lag_rsp_ff), fabric_lag.prev_control_state_0);
  mkConnection(toClient(fwd_result_req_ff, fwd_result_rsp_ff), fwd_result.prev_control_state_0);
  mkConnection(toClient(ingress_bd_stats_req_ff, ingress_bd_stats_rsp_ff), ingress_bd_stats.prev_control_state_0);
  mkConnection(toClient(ingress_port_mapping_req_ff, ingress_port_mapping_rsp_ff), ingress_port_mapping.prev_control_state_0);
  mkConnection(toClient(ingress_port_properties_req_ff, ingress_port_properties_rsp_ff), ingress_port_properties.prev_control_state_0);
  mkConnection(toClient(int_sink_update_outer_req_ff, int_sink_update_outer_rsp_ff), int_sink_update_outer.prev_control_state_0);
  mkConnection(toClient(int_source_req_ff, int_source_rsp_ff), int_source.prev_control_state_0);
  mkConnection(toClient(int_terminate_req_ff, int_terminate_rsp_ff), int_terminate.prev_control_state_0);
  mkConnection(toClient(ip_acl_req_ff, ip_acl_rsp_ff), ip_acl.prev_control_state_0);
  mkConnection(toClient(ipsg_req_ff, ipsg_rsp_ff), ipsg.prev_control_state_0);
  mkConnection(toClient(ipsg_permit_special_req_ff, ipsg_permit_special_rsp_ff), ipsg_permit_special.prev_control_state_0);
  mkConnection(toClient(ipv4_dest_vtep_req_ff, ipv4_dest_vtep_rsp_ff), ipv4_dest_vtep.prev_control_state_0);
  mkConnection(toClient(ipv4_fib_req_ff, ipv4_fib_rsp_ff), ipv4_fib.prev_control_state_0);
  mkConnection(toClient(ipv4_fib_lpm_req_ff, ipv4_fib_lpm_rsp_ff), ipv4_fib_lpm.prev_control_state_0);
  mkConnection(toClient(ipv4_multicast_bridge_req_ff, ipv4_multicast_bridge_rsp_ff), ipv4_multicast_bridge.prev_control_state_0);
  mkConnection(toClient(ipv4_multicast_bridge_star_g_req_ff, ipv4_multicast_bridge_star_g_rsp_ff), ipv4_multicast_bridge_star_g.prev_control_state_0);
  mkConnection(toClient(ipv4_multicast_route_req_ff, ipv4_multicast_route_rsp_ff), ipv4_multicast_route.prev_control_state_0);
  mkConnection(toClient(ipv4_multicast_route_star_g_req_ff, ipv4_multicast_route_star_g_rsp_ff), ipv4_multicast_route_star_g.prev_control_state_0);
  mkConnection(toClient(ipv4_racl_req_ff, ipv4_racl_rsp_ff), ipv4_racl.prev_control_state_0);
  mkConnection(toClient(ipv4_src_vtep_req_ff, ipv4_src_vtep_rsp_ff), ipv4_src_vtep.prev_control_state_0);
  mkConnection(toClient(ipv4_urpf_req_ff, ipv4_urpf_rsp_ff), ipv4_urpf.prev_control_state_0);
  mkConnection(toClient(ipv4_urpf_lpm_req_ff, ipv4_urpf_lpm_rsp_ff), ipv4_urpf_lpm.prev_control_state_0);
  mkConnection(toClient(ipv6_acl_req_ff, ipv6_acl_rsp_ff), ipv6_acl.prev_control_state_0);
  mkConnection(toClient(ipv6_dest_vtep_req_ff, ipv6_dest_vtep_rsp_ff), ipv6_dest_vtep.prev_control_state_0);
  mkConnection(toClient(ipv6_fib_req_ff, ipv6_fib_rsp_ff), ipv6_fib.prev_control_state_0);
  mkConnection(toClient(ipv6_fib_lpm_req_ff, ipv6_fib_lpm_rsp_ff), ipv6_fib_lpm.prev_control_state_0);
  mkConnection(toClient(ipv6_multicast_bridge_req_ff, ipv6_multicast_bridge_rsp_ff), ipv6_multicast_bridge.prev_control_state_0);
  mkConnection(toClient(ipv6_multicast_bridge_star_g_req_ff, ipv6_multicast_bridge_star_g_rsp_ff), ipv6_multicast_bridge_star_g.prev_control_state_0);
  mkConnection(toClient(ipv6_multicast_route_req_ff, ipv6_multicast_route_rsp_ff), ipv6_multicast_route.prev_control_state_0);
  mkConnection(toClient(ipv6_multicast_route_star_g_req_ff, ipv6_multicast_route_star_g_rsp_ff), ipv6_multicast_route_star_g.prev_control_state_0);
  mkConnection(toClient(ipv6_racl_req_ff, ipv6_racl_rsp_ff), ipv6_racl.prev_control_state_0);
  mkConnection(toClient(ipv6_src_vtep_req_ff, ipv6_src_vtep_rsp_ff), ipv6_src_vtep.prev_control_state_0);
  mkConnection(toClient(ipv6_urpf_req_ff, ipv6_urpf_rsp_ff), ipv6_urpf.prev_control_state_0);
  mkConnection(toClient(ipv6_urpf_lpm_req_ff, ipv6_urpf_lpm_rsp_ff), ipv6_urpf_lpm.prev_control_state_0);
  mkConnection(toClient(lag_group_req_ff, lag_group_rsp_ff), lag_group.prev_control_state_0);
  mkConnection(toClient(learn_notify_req_ff, learn_notify_rsp_ff), learn_notify.prev_control_state_0);
  mkConnection(toClient(mac_acl_req_ff, mac_acl_rsp_ff), mac_acl.prev_control_state_0);
  mkConnection(toClient(meter_action_req_ff, meter_action_rsp_ff), meter_action.prev_control_state_0);
  mkConnection(toClient(meter_index_req_ff, meter_index_rsp_ff), meter_index.prev_control_state_0);
  mkConnection(toClient(mpls_req_ff, mpls_rsp_ff), mpls.prev_control_state_0);
  mkConnection(toClient(native_packet_over_fabric_req_ff, native_packet_over_fabric_rsp_ff), native_packet_over_fabric.prev_control_state_0);
  mkConnection(toClient(nexthop_req_ff, nexthop_rsp_ff), nexthop.prev_control_state_0);
  mkConnection(toClient(outer_ipv4_multicast_req_ff, outer_ipv4_multicast_rsp_ff), outer_ipv4_multicast.prev_control_state_0);
  mkConnection(toClient(outer_ipv4_multicast_star_g_req_ff, outer_ipv4_multicast_star_g_rsp_ff), outer_ipv4_multicast_star_g.prev_control_state_0);
  mkConnection(toClient(outer_ipv6_multicast_req_ff, outer_ipv6_multicast_rsp_ff), outer_ipv6_multicast.prev_control_state_0);
  mkConnection(toClient(outer_ipv6_multicast_star_g_req_ff, outer_ipv6_multicast_star_g_rsp_ff), outer_ipv6_multicast_star_g.prev_control_state_0);
  mkConnection(toClient(outer_rmac_req_ff, outer_rmac_rsp_ff), outer_rmac.prev_control_state_0);
  mkConnection(toClient(port_vlan_mapping_req_ff, port_vlan_mapping_rsp_ff), port_vlan_mapping.prev_control_state_0);
  mkConnection(toClient(qos_req_ff, qos_rsp_ff), qos.prev_control_state_0);
  mkConnection(toClient(rmac_req_ff, rmac_rsp_ff), rmac.prev_control_state_0);
  mkConnection(toClient(sflow_ing_take_sample_req_ff, sflow_ing_take_sample_rsp_ff), sflow_ing_take_sample.prev_control_state_0);
  mkConnection(toClient(sflow_ingress_req_ff, sflow_ingress_rsp_ff), sflow_ingress.prev_control_state_0);
  mkConnection(toClient(smac_req_ff, smac_rsp_ff), smac.prev_control_state_0);
  mkConnection(toClient(spanning_tree_req_ff, spanning_tree_rsp_ff), spanning_tree.prev_control_state_0);
  mkConnection(toClient(storm_control_req_ff, storm_control_rsp_ff), storm_control.prev_control_state_0);
  mkConnection(toClient(storm_control_stats_req_ff, storm_control_stats_rsp_ff), storm_control_stats.prev_control_state_0);
  mkConnection(toClient(switch_config_params_req_ff, switch_config_params_rsp_ff), switch_config_params.prev_control_state_0);
  mkConnection(toClient(system_acl_req_ff, system_acl_rsp_ff), system_acl.prev_control_state_0);
  mkConnection(toClient(tunnel_req_ff, tunnel_rsp_ff), tunnel.prev_control_state_0);
  mkConnection(toClient(tunnel_lookup_miss_req_ff, tunnel_lookup_miss_rsp_ff), tunnel_lookup_miss.prev_control_state_0);
  mkConnection(toClient(tunnel_miss_req_ff, tunnel_miss_rsp_ff), tunnel_miss.prev_control_state_0);
  mkConnection(toClient(urpf_bd_req_ff, urpf_bd_rsp_ff), urpf_bd.prev_control_state_0);
  mkConnection(toClient(validate_mpls_packet_req_ff, validate_mpls_packet_rsp_ff), validate_mpls_packet.prev_control_state_0);
  mkConnection(toClient(validate_outer_ethernet_req_ff, validate_outer_ethernet_rsp_ff), validate_outer_ethernet.prev_control_state_0);
  mkConnection(toClient(validate_outer_ipv4_packet_req_ff, validate_outer_ipv4_packet_rsp_ff), validate_outer_ipv4_packet.prev_control_state_0);
  mkConnection(toClient(validate_outer_ipv6_packet_req_ff, validate_outer_ipv6_packet_rsp_ff), validate_outer_ipv6_packet.prev_control_state_0);
  mkConnection(toClient(validate_packet_req_ff, validate_packet_rsp_ff), validate_packet.prev_control_state_0);
  // Basic Blocks
  AclStatsUpdate acl_stats_update_0 <- mkAclStatsUpdate();
  Nop nop_0 <- mkNop();
  SetBdFloodMcIndex set_bd_flood_mc_index_0 <- mkSetBdFloodMcIndex();
  ComputeLkpIpv4Hash compute_lkp_ipv4_hash_0 <- mkComputeLkpIpv4Hash();
  ComputeLkpIpv6Hash compute_lkp_ipv6_hash_0 <- mkComputeLkpIpv6Hash();
  ComputeLkpNonIpHash compute_lkp_non_ip_hash_0 <- mkComputeLkpNonIpHash();
  ComputedTwoHashes computed_two_hashes_0 <- mkComputedTwoHashes();
  ComputedOneHash computed_one_hash_0 <- mkComputedOneHash();
  Nop nop_1 <- mkNop();
  DmacHit dmac_hit_0 <- mkDmacHit();
  DmacMulticastHit dmac_multicast_hit_0 <- mkDmacMulticastHit();
  DmacMiss dmac_miss_0 <- mkDmacMiss();
  DmacRedirectNexthop dmac_redirect_nexthop_0 <- mkDmacRedirectNexthop();
  DmacRedirectEcmp dmac_redirect_ecmp_0 <- mkDmacRedirectEcmp();
  DmacDrop dmac_drop_0 <- mkDmacDrop();
  DropStatsUpdate drop_stats_update_0 <- mkDropStatsUpdate();
  Nop nop_2 <- mkNop();
  SetEcmpNexthopDetails set_ecmp_nexthop_details_0 <- mkSetEcmpNexthopDetails();
  SetEcmpNexthopDetailsForPostRoutedFlood set_ecmp_nexthop_details_for_post_routed_flood_0 <- mkSetEcmpNexthopDetailsForPostRoutedFlood();
  Nop nop_3 <- mkNop();
  TerminateCpuPacket terminate_cpu_packet_0 <- mkTerminateCpuPacket();
  SwitchFabricUnicastPacket switch_fabric_unicast_packet_0 <- mkSwitchFabricUnicastPacket();
  TerminateFabricUnicastPacket terminate_fabric_unicast_packet_0 <- mkTerminateFabricUnicastPacket();
  SwitchFabricMulticastPacket switch_fabric_multicast_packet_0 <- mkSwitchFabricMulticastPacket();
  TerminateFabricMulticastPacket terminate_fabric_multicast_packet_0 <- mkTerminateFabricMulticastPacket();
  Nop nop_4 <- mkNop();
  SetIngressIfindexProperties set_ingress_ifindex_properties_0 <- mkSetIngressIfindexProperties();
  Nop nop_5 <- mkNop();
  SetFabricLagPort set_fabric_lag_port_0 <- mkSetFabricLagPort();
  SetFabricMulticast set_fabric_multicast_0 <- mkSetFabricMulticast();
  Nop nop_6 <- mkNop();
  SetL2RedirectAction set_l2_redirect_action_0 <- mkSetL2RedirectAction();
  SetFibRedirectAction set_fib_redirect_action_0 <- mkSetFibRedirectAction();
  SetCpuRedirectAction set_cpu_redirect_action_0 <- mkSetCpuRedirectAction();
  SetAclRedirectAction set_acl_redirect_action_0 <- mkSetAclRedirectAction();
  SetRaclRedirectAction set_racl_redirect_action_0 <- mkSetRaclRedirectAction();
  SetMulticastRouteAction set_multicast_route_action_0 <- mkSetMulticastRouteAction();
  SetMulticastBridgeAction set_multicast_bridge_action_0 <- mkSetMulticastBridgeAction();
  SetMulticastFlood set_multicast_flood_0 <- mkSetMulticastFlood();
  SetMulticastDrop set_multicast_drop_0 <- mkSetMulticastDrop();
  UpdateIngressBdStats update_ingress_bd_stats_0 <- mkUpdateIngressBdStats();
  SetIfindex set_ifindex_0 <- mkSetIfindex();
  SetIngressPortProperties set_ingress_port_properties_0 <- mkSetIngressPortProperties();
  IntSinkUpdateVxlanGpeV4 int_sink_update_vxlan_gpe_v4_0 <- mkIntSinkUpdateVxlanGpeV4();
  Nop nop_7 <- mkNop();
  IntSetSrc int_set_src_0 <- mkIntSetSrc();
  IntSetNoSrc int_set_no_src_0 <- mkIntSetNoSrc();
  IntSinkGpe int_sink_gpe_0 <- mkIntSinkGpe();
  IntNoSink int_no_sink_0 <- mkIntNoSink();
  Nop nop_8 <- mkNop();
  AclDeny acl_deny_0 <- mkAclDeny();
  AclPermit acl_permit_0 <- mkAclPermit();
  AclMirror acl_mirror_0 <- mkAclMirror();
  AclRedirectNexthop acl_redirect_nexthop_0 <- mkAclRedirectNexthop();
  AclRedirectEcmp acl_redirect_ecmp_0 <- mkAclRedirectEcmp();
  OnMiss on_miss_0 <- mkOnMiss();
  IpsgMiss ipsg_miss_0 <- mkIpsgMiss();
  Nop nop_9 <- mkNop();
  SetTunnelTerminationFlag set_tunnel_termination_flag_0 <- mkSetTunnelTerminationFlag();
  SetTunnelVniAndTerminationFlag set_tunnel_vni_and_termination_flag_0 <- mkSetTunnelVniAndTerminationFlag();
  OnMiss on_miss_1 <- mkOnMiss();
  FibHitNexthop fib_hit_nexthop_0 <- mkFibHitNexthop();
  FibHitEcmp fib_hit_ecmp_0 <- mkFibHitEcmp();
  OnMiss on_miss_2 <- mkOnMiss();
  FibHitNexthop fib_hit_nexthop_1 <- mkFibHitNexthop();
  FibHitEcmp fib_hit_ecmp_1 <- mkFibHitEcmp();
  OnMiss on_miss_3 <- mkOnMiss();
  MulticastBridgeSGHit multicast_bridge_s_g_hit_0 <- mkMulticastBridgeSGHit();
  Nop nop_10 <- mkNop();
  MulticastBridgeStarGHit multicast_bridge_star_g_hit_0 <- mkMulticastBridgeStarGHit();
  OnMiss on_miss_4 <- mkOnMiss();
  MulticastRouteSGHit multicast_route_s_g_hit_0 <- mkMulticastRouteSGHit();
  MulticastRouteStarGMiss multicast_route_star_g_miss_0 <- mkMulticastRouteStarGMiss();
  MulticastRouteSmStarGHit multicast_route_sm_star_g_hit_0 <- mkMulticastRouteSmStarGHit();
  MulticastRouteBidirStarGHit multicast_route_bidir_star_g_hit_0 <- mkMulticastRouteBidirStarGHit();
  Nop nop_11 <- mkNop();
  RaclDeny racl_deny_0 <- mkRaclDeny();
  RaclPermit racl_permit_0 <- mkRaclPermit();
  RaclRedirectNexthop racl_redirect_nexthop_0 <- mkRaclRedirectNexthop();
  RaclRedirectEcmp racl_redirect_ecmp_0 <- mkRaclRedirectEcmp();
  OnMiss on_miss_5 <- mkOnMiss();
  SrcVtepHit src_vtep_hit_0 <- mkSrcVtepHit();
  OnMiss on_miss_6 <- mkOnMiss();
  Ipv4UrpfHit ipv4_urpf_hit_0 <- mkIpv4UrpfHit();
  Ipv4UrpfHit ipv4_urpf_hit_1 <- mkIpv4UrpfHit();
  UrpfMiss urpf_miss_0 <- mkUrpfMiss();
  Nop nop_12 <- mkNop();
  AclDeny acl_deny_1 <- mkAclDeny();
  AclPermit acl_permit_1 <- mkAclPermit();
  AclMirror acl_mirror_1 <- mkAclMirror();
  AclRedirectNexthop acl_redirect_nexthop_1 <- mkAclRedirectNexthop();
  AclRedirectEcmp acl_redirect_ecmp_1 <- mkAclRedirectEcmp();
  Nop nop_13 <- mkNop();
  SetTunnelTerminationFlag set_tunnel_termination_flag_1 <- mkSetTunnelTerminationFlag();
  SetTunnelVniAndTerminationFlag set_tunnel_vni_and_termination_flag_1 <- mkSetTunnelVniAndTerminationFlag();
  OnMiss on_miss_7 <- mkOnMiss();
  FibHitNexthop fib_hit_nexthop_2 <- mkFibHitNexthop();
  FibHitEcmp fib_hit_ecmp_2 <- mkFibHitEcmp();
  OnMiss on_miss_8 <- mkOnMiss();
  FibHitNexthop fib_hit_nexthop_3 <- mkFibHitNexthop();
  FibHitEcmp fib_hit_ecmp_3 <- mkFibHitEcmp();
  OnMiss on_miss_9 <- mkOnMiss();
  MulticastBridgeSGHit multicast_bridge_s_g_hit_1 <- mkMulticastBridgeSGHit();
  Nop nop_14 <- mkNop();
  MulticastBridgeStarGHit multicast_bridge_star_g_hit_1 <- mkMulticastBridgeStarGHit();
  OnMiss on_miss_10 <- mkOnMiss();
  MulticastRouteSGHit multicast_route_s_g_hit_1 <- mkMulticastRouteSGHit();
  MulticastRouteStarGMiss multicast_route_star_g_miss_1 <- mkMulticastRouteStarGMiss();
  MulticastRouteSmStarGHit multicast_route_sm_star_g_hit_1 <- mkMulticastRouteSmStarGHit();
  MulticastRouteBidirStarGHit multicast_route_bidir_star_g_hit_1 <- mkMulticastRouteBidirStarGHit();
  Nop nop_15 <- mkNop();
  RaclDeny racl_deny_1 <- mkRaclDeny();
  RaclPermit racl_permit_1 <- mkRaclPermit();
  RaclRedirectNexthop racl_redirect_nexthop_1 <- mkRaclRedirectNexthop();
  RaclRedirectEcmp racl_redirect_ecmp_1 <- mkRaclRedirectEcmp();
  OnMiss on_miss_11 <- mkOnMiss();
  SrcVtepHit src_vtep_hit_1 <- mkSrcVtepHit();
  OnMiss on_miss_12 <- mkOnMiss();
  Ipv6UrpfHit ipv6_urpf_hit_0 <- mkIpv6UrpfHit();
  Ipv6UrpfHit ipv6_urpf_hit_1 <- mkIpv6UrpfHit();
  UrpfMiss urpf_miss_1 <- mkUrpfMiss();
  SetLagMiss set_lag_miss_0 <- mkSetLagMiss();
  SetLagPort set_lag_port_0 <- mkSetLagPort();
  SetLagRemotePort set_lag_remote_port_0 <- mkSetLagRemotePort();
  Nop nop_16 <- mkNop();
  GenerateLearnNotify generate_learn_notify_0 <- mkGenerateLearnNotify();
  Nop nop_17 <- mkNop();
  AclDeny acl_deny_2 <- mkAclDeny();
  AclPermit acl_permit_2 <- mkAclPermit();
  AclMirror acl_mirror_2 <- mkAclMirror();
  AclRedirectNexthop acl_redirect_nexthop_2 <- mkAclRedirectNexthop();
  AclRedirectEcmp acl_redirect_ecmp_2 <- mkAclRedirectEcmp();
  MeterPermit meter_permit_0 <- mkMeterPermit();
  MeterDeny meter_deny_0 <- mkMeterDeny();
  Nop nop_18 <- mkNop();
  TerminateEompls terminate_eompls_0 <- mkTerminateEompls();
  TerminateVpls terminate_vpls_0 <- mkTerminateVpls();
  TerminateIpv4OverMpls terminate_ipv4_over_mpls_0 <- mkTerminateIpv4OverMpls();
  TerminateIpv6OverMpls terminate_ipv6_over_mpls_0 <- mkTerminateIpv6OverMpls();
  TerminatePw terminate_pw_0 <- mkTerminatePw();
  ForwardMpls forward_mpls_0 <- mkForwardMpls();
  NonIpOverFabric non_ip_over_fabric_0 <- mkNonIpOverFabric();
  Ipv4OverFabric ipv4_over_fabric_0 <- mkIpv4OverFabric();
  Ipv6OverFabric ipv6_over_fabric_0 <- mkIpv6OverFabric();
  Nop nop_19 <- mkNop();
  SetNexthopDetails set_nexthop_details_0 <- mkSetNexthopDetails();
  SetNexthopDetailsForPostRoutedFlood set_nexthop_details_for_post_routed_flood_0 <- mkSetNexthopDetailsForPostRoutedFlood();
  Nop nop_20 <- mkNop();
  OnMiss on_miss_13 <- mkOnMiss();
  OuterMulticastRouteSGHit outer_multicast_route_s_g_hit_0 <- mkOuterMulticastRouteSGHit();
  OuterMulticastBridgeSGHit outer_multicast_bridge_s_g_hit_0 <- mkOuterMulticastBridgeSGHit();
  Nop nop_21 <- mkNop();
  OuterMulticastRouteSmStarGHit outer_multicast_route_sm_star_g_hit_0 <- mkOuterMulticastRouteSmStarGHit();
  OuterMulticastRouteBidirStarGHit outer_multicast_route_bidir_star_g_hit_0 <- mkOuterMulticastRouteBidirStarGHit();
  OuterMulticastBridgeStarGHit outer_multicast_bridge_star_g_hit_0 <- mkOuterMulticastBridgeStarGHit();
  Nop nop_22 <- mkNop();
  OnMiss on_miss_14 <- mkOnMiss();
  OuterMulticastRouteSGHit outer_multicast_route_s_g_hit_1 <- mkOuterMulticastRouteSGHit();
  OuterMulticastBridgeSGHit outer_multicast_bridge_s_g_hit_1 <- mkOuterMulticastBridgeSGHit();
  Nop nop_23 <- mkNop();
  OuterMulticastRouteSmStarGHit outer_multicast_route_sm_star_g_hit_1 <- mkOuterMulticastRouteSmStarGHit();
  OuterMulticastRouteBidirStarGHit outer_multicast_route_bidir_star_g_hit_1 <- mkOuterMulticastRouteBidirStarGHit();
  OuterMulticastBridgeStarGHit outer_multicast_bridge_star_g_hit_1 <- mkOuterMulticastBridgeStarGHit();
  OnMiss on_miss_15 <- mkOnMiss();
  OuterRmacHit outer_rmac_hit_0 <- mkOuterRmacHit();
  SetBdProperties set_bd_properties_0 <- mkSetBdProperties();
  PortVlanMappingMiss port_vlan_mapping_miss_0 <- mkPortVlanMappingMiss();
  Nop nop_24 <- mkNop();
  ApplyCosMarking apply_cos_marking_0 <- mkApplyCosMarking();
  ApplyDscpMarking apply_dscp_marking_0 <- mkApplyDscpMarking();
  ApplyTcMarking apply_tc_marking_0 <- mkApplyTcMarking();
  RmacHit rmac_hit_0 <- mkRmacHit();
  RmacMiss rmac_miss_0 <- mkRmacMiss();
  Nop nop_25 <- mkNop();
  SflowIngPktToCpu sflow_ing_pkt_to_cpu_0 <- mkSflowIngPktToCpu();
  Nop nop_26 <- mkNop();
  SflowIngSessionEnable sflow_ing_session_enable_0 <- mkSflowIngSessionEnable();
  Nop nop_27 <- mkNop();
  SmacMiss smac_miss_0 <- mkSmacMiss();
  SmacHit smac_hit_0 <- mkSmacHit();
  SetStpState set_stp_state_0 <- mkSetStpState();
  Nop nop_28 <- mkNop();
  SetStormControlMeter set_storm_control_meter_0 <- mkSetStormControlMeter();
  Nop nop_29 <- mkNop();
  SetConfigParameters set_config_parameters_0 <- mkSetConfigParameters();
  Nop nop_30 <- mkNop();
  RedirectToCpu redirect_to_cpu_0 <- mkRedirectToCpu();
  CopyToCpuWithReason copy_to_cpu_with_reason_0 <- mkCopyToCpuWithReason();
  CopyToCpu copy_to_cpu_0 <- mkCopyToCpu();
  DropPacket drop_packet_0 <- mkDropPacket();
  DropPacketWithReason drop_packet_with_reason_0 <- mkDropPacketWithReason();
  NegativeMirror negative_mirror_0 <- mkNegativeMirror();
  Nop nop_31 <- mkNop();
  ATunnelLookupMiss tunnel_lookup_miss_0 <- mkATunnelLookupMiss();
  TerminateTunnelInnerNonIp terminate_tunnel_inner_non_ip_0 <- mkTerminateTunnelInnerNonIp();
  TerminateTunnelInnerEthernetIpv4 terminate_tunnel_inner_ethernet_ipv4_0 <- mkTerminateTunnelInnerEthernetIpv4();
  TerminateTunnelInnerIpv4 terminate_tunnel_inner_ipv4_0 <- mkTerminateTunnelInnerIpv4();
  TerminateTunnelInnerEthernetIpv6 terminate_tunnel_inner_ethernet_ipv6_0 <- mkTerminateTunnelInnerEthernetIpv6();
  TerminateTunnelInnerIpv6 terminate_tunnel_inner_ipv6_0 <- mkTerminateTunnelInnerIpv6();
  NonIpTunnelLookupMiss non_ip_tunnel_lookup_miss_0 <- mkNonIpTunnelLookupMiss();
  Ipv4TunnelLookupMiss ipv4_tunnel_lookup_miss_0 <- mkIpv4TunnelLookupMiss();
  Ipv6TunnelLookupMiss ipv6_tunnel_lookup_miss_0 <- mkIpv6TunnelLookupMiss();
  NonIpTunnelLookupMiss non_ip_tunnel_lookup_miss_1 <- mkNonIpTunnelLookupMiss();
  Ipv4TunnelLookupMiss ipv4_tunnel_lookup_miss_1 <- mkIpv4TunnelLookupMiss();
  Ipv6TunnelLookupMiss ipv6_tunnel_lookup_miss_1 <- mkIpv6TunnelLookupMiss();
  Nop nop_32 <- mkNop();
  UrpfBdMiss urpf_bd_miss_0 <- mkUrpfBdMiss();
  SetValidMplsLabel1 set_valid_mpls_label1_0 <- mkSetValidMplsLabel1();
  SetValidMplsLabel2 set_valid_mpls_label2_0 <- mkSetValidMplsLabel2();
  SetValidMplsLabel3 set_valid_mpls_label3_0 <- mkSetValidMplsLabel3();
  MalformedOuterEthernetPacket malformed_outer_ethernet_packet_0 <- mkMalformedOuterEthernetPacket();
  SetValidOuterUnicastPacketUntagged set_valid_outer_unicast_packet_untagged_0 <- mkSetValidOuterUnicastPacketUntagged();
  SetValidOuterUnicastPacketSingleTagged set_valid_outer_unicast_packet_single_tagged_0 <- mkSetValidOuterUnicastPacketSingleTagged();
  SetValidOuterUnicastPacketDoubleTagged set_valid_outer_unicast_packet_double_tagged_0 <- mkSetValidOuterUnicastPacketDoubleTagged();
  SetValidOuterUnicastPacketQinqTagged set_valid_outer_unicast_packet_qinq_tagged_0 <- mkSetValidOuterUnicastPacketQinqTagged();
  SetValidOuterMulticastPacketUntagged set_valid_outer_multicast_packet_untagged_0 <- mkSetValidOuterMulticastPacketUntagged();
  SetValidOuterMulticastPacketSingleTagged set_valid_outer_multicast_packet_single_tagged_0 <- mkSetValidOuterMulticastPacketSingleTagged();
  SetValidOuterMulticastPacketDoubleTagged set_valid_outer_multicast_packet_double_tagged_0 <- mkSetValidOuterMulticastPacketDoubleTagged();
  SetValidOuterMulticastPacketQinqTagged set_valid_outer_multicast_packet_qinq_tagged_0 <- mkSetValidOuterMulticastPacketQinqTagged();
  SetValidOuterBroadcastPacketUntagged set_valid_outer_broadcast_packet_untagged_0 <- mkSetValidOuterBroadcastPacketUntagged();
  SetValidOuterBroadcastPacketSingleTagged set_valid_outer_broadcast_packet_single_tagged_0 <- mkSetValidOuterBroadcastPacketSingleTagged();
  SetValidOuterBroadcastPacketDoubleTagged set_valid_outer_broadcast_packet_double_tagged_0 <- mkSetValidOuterBroadcastPacketDoubleTagged();
  SetValidOuterBroadcastPacketQinqTagged set_valid_outer_broadcast_packet_qinq_tagged_0 <- mkSetValidOuterBroadcastPacketQinqTagged();
  SetValidOuterIpv4Packet set_valid_outer_ipv4_packet_0 <- mkSetValidOuterIpv4Packet();
  SetMalformedOuterIpv4Packet set_malformed_outer_ipv4_packet_0 <- mkSetMalformedOuterIpv4Packet();
  SetValidOuterIpv6Packet set_valid_outer_ipv6_packet_0 <- mkSetValidOuterIpv6Packet();
  SetMalformedOuterIpv6Packet set_malformed_outer_ipv6_packet_0 <- mkSetMalformedOuterIpv6Packet();
  Nop nop_33 <- mkNop();
  SetUnicast set_unicast_0 <- mkSetUnicast();
  SetUnicastAndIpv6SrcIsLinkLocal set_unicast_and_ipv6_src_is_link_local_0 <- mkSetUnicastAndIpv6SrcIsLinkLocal();
  SetMulticast set_multicast_0 <- mkSetMulticast();
  SetMulticastAndIpv6SrcIsLinkLocal set_multicast_and_ipv6_src_is_link_local_0 <- mkSetMulticastAndIpv6SrcIsLinkLocal();
  SetBroadcast set_broadcast_0 <- mkSetBroadcast();
  SetMalformedPacket set_malformed_packet_0 <- mkSetMalformedPacket();
  mkChan(mkFIFOF, mkFIFOF, acl_stats.next_control_state_0, acl_stats_update_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, bd_flood.next_control_state_0, nop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, bd_flood.next_control_state_1, set_bd_flood_mc_index_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, compute_ipv4_hashes.next_control_state_0, compute_lkp_ipv4_hash_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, compute_ipv6_hashes.next_control_state_0, compute_lkp_ipv6_hash_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, compute_non_ip_hashes.next_control_state_0, compute_lkp_non_ip_hash_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, compute_other_hashes.next_control_state_0, computed_two_hashes_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, compute_other_hashes.next_control_state_1, computed_one_hash_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, dmac.next_control_state_0, nop_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, dmac.next_control_state_1, dmac_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, dmac.next_control_state_2, dmac_multicast_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, dmac.next_control_state_3, dmac_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, dmac.next_control_state_4, dmac_redirect_nexthop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, dmac.next_control_state_5, dmac_redirect_ecmp_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, dmac.next_control_state_6, dmac_drop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, drop_stats.next_control_state_0, drop_stats_update_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ecmp_group.next_control_state_0, nop_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ecmp_group.next_control_state_1, set_ecmp_nexthop_details_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ecmp_group.next_control_state_2, set_ecmp_nexthop_details_for_post_routed_flood_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_ingress_dst_lkp.next_control_state_0, nop_3.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_ingress_dst_lkp.next_control_state_1, terminate_cpu_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_ingress_dst_lkp.next_control_state_2, switch_fabric_unicast_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_ingress_dst_lkp.next_control_state_3, terminate_fabric_unicast_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_ingress_dst_lkp.next_control_state_4, switch_fabric_multicast_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_ingress_dst_lkp.next_control_state_5, terminate_fabric_multicast_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_ingress_src_lkp.next_control_state_0, nop_4.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_ingress_src_lkp.next_control_state_1, set_ingress_ifindex_properties_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_lag.next_control_state_0, nop_5.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_lag.next_control_state_1, set_fabric_lag_port_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fabric_lag.next_control_state_2, set_fabric_multicast_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_0, nop_6.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_1, set_l2_redirect_action_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_2, set_fib_redirect_action_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_3, set_cpu_redirect_action_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_4, set_acl_redirect_action_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_5, set_racl_redirect_action_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_6, set_multicast_route_action_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_7, set_multicast_bridge_action_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_8, set_multicast_flood_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, fwd_result.next_control_state_9, set_multicast_drop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ingress_bd_stats.next_control_state_0, update_ingress_bd_stats_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ingress_port_mapping.next_control_state_0, set_ifindex_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ingress_port_properties.next_control_state_0, set_ingress_port_properties_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_sink_update_outer.next_control_state_0, int_sink_update_vxlan_gpe_v4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_sink_update_outer.next_control_state_1, nop_7.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_source.next_control_state_0, int_set_src_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_source.next_control_state_1, int_set_no_src_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_terminate.next_control_state_0, int_sink_gpe_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_terminate.next_control_state_1, int_no_sink_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ip_acl.next_control_state_0, nop_8.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ip_acl.next_control_state_1, acl_deny_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ip_acl.next_control_state_2, acl_permit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ip_acl.next_control_state_3, acl_mirror_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ip_acl.next_control_state_4, acl_redirect_nexthop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ip_acl.next_control_state_5, acl_redirect_ecmp_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipsg.next_control_state_0, on_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipsg_permit_special.next_control_state_0, ipsg_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_dest_vtep.next_control_state_0, nop_9.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_dest_vtep.next_control_state_1, set_tunnel_termination_flag_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_dest_vtep.next_control_state_2, set_tunnel_vni_and_termination_flag_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_fib.next_control_state_0, on_miss_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_fib.next_control_state_1, fib_hit_nexthop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_fib.next_control_state_2, fib_hit_ecmp_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_fib_lpm.next_control_state_0, on_miss_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_fib_lpm.next_control_state_1, fib_hit_nexthop_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_fib_lpm.next_control_state_2, fib_hit_ecmp_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_bridge.next_control_state_0, on_miss_3.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_bridge.next_control_state_1, multicast_bridge_s_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_bridge_star_g.next_control_state_0, nop_10.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_bridge_star_g.next_control_state_1, multicast_bridge_star_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_route.next_control_state_0, on_miss_4.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_route.next_control_state_1, multicast_route_s_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_route_star_g.next_control_state_0, multicast_route_star_g_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_route_star_g.next_control_state_1, multicast_route_sm_star_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_multicast_route_star_g.next_control_state_2, multicast_route_bidir_star_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_racl.next_control_state_0, nop_11.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_racl.next_control_state_1, racl_deny_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_racl.next_control_state_2, racl_permit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_racl.next_control_state_3, racl_redirect_nexthop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_racl.next_control_state_4, racl_redirect_ecmp_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_src_vtep.next_control_state_0, on_miss_5.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_src_vtep.next_control_state_1, src_vtep_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_urpf.next_control_state_0, on_miss_6.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_urpf.next_control_state_1, ipv4_urpf_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_urpf_lpm.next_control_state_0, ipv4_urpf_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv4_urpf_lpm.next_control_state_1, urpf_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_acl.next_control_state_0, nop_12.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_acl.next_control_state_1, acl_deny_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_acl.next_control_state_2, acl_permit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_acl.next_control_state_3, acl_mirror_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_acl.next_control_state_4, acl_redirect_nexthop_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_acl.next_control_state_5, acl_redirect_ecmp_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_dest_vtep.next_control_state_0, nop_13.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_dest_vtep.next_control_state_1, set_tunnel_termination_flag_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_dest_vtep.next_control_state_2, set_tunnel_vni_and_termination_flag_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_fib.next_control_state_0, on_miss_7.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_fib.next_control_state_1, fib_hit_nexthop_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_fib.next_control_state_2, fib_hit_ecmp_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_fib_lpm.next_control_state_0, on_miss_8.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_fib_lpm.next_control_state_1, fib_hit_nexthop_3.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_fib_lpm.next_control_state_2, fib_hit_ecmp_3.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_bridge.next_control_state_0, on_miss_9.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_bridge.next_control_state_1, multicast_bridge_s_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_bridge_star_g.next_control_state_0, nop_14.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_bridge_star_g.next_control_state_1, multicast_bridge_star_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_route.next_control_state_0, on_miss_10.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_route.next_control_state_1, multicast_route_s_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_route_star_g.next_control_state_0, multicast_route_star_g_miss_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_route_star_g.next_control_state_1, multicast_route_sm_star_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_multicast_route_star_g.next_control_state_2, multicast_route_bidir_star_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_racl.next_control_state_0, nop_15.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_racl.next_control_state_1, racl_deny_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_racl.next_control_state_2, racl_permit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_racl.next_control_state_3, racl_redirect_nexthop_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_racl.next_control_state_4, racl_redirect_ecmp_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_src_vtep.next_control_state_0, on_miss_11.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_src_vtep.next_control_state_1, src_vtep_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_urpf.next_control_state_0, on_miss_12.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_urpf.next_control_state_1, ipv6_urpf_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_urpf_lpm.next_control_state_0, ipv6_urpf_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, ipv6_urpf_lpm.next_control_state_1, urpf_miss_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, lag_group.next_control_state_0, set_lag_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, lag_group.next_control_state_1, set_lag_port_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, lag_group.next_control_state_2, set_lag_remote_port_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, learn_notify.next_control_state_0, nop_16.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, learn_notify.next_control_state_1, generate_learn_notify_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mac_acl.next_control_state_0, nop_17.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mac_acl.next_control_state_1, acl_deny_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mac_acl.next_control_state_2, acl_permit_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mac_acl.next_control_state_3, acl_mirror_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mac_acl.next_control_state_4, acl_redirect_nexthop_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mac_acl.next_control_state_5, acl_redirect_ecmp_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, meter_action.next_control_state_0, meter_permit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, meter_action.next_control_state_1, meter_deny_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, meter_index.next_control_state_0, nop_18.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mpls.next_control_state_0, terminate_eompls_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mpls.next_control_state_1, terminate_vpls_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mpls.next_control_state_2, terminate_ipv4_over_mpls_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mpls.next_control_state_3, terminate_ipv6_over_mpls_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mpls.next_control_state_4, terminate_pw_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mpls.next_control_state_5, forward_mpls_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, native_packet_over_fabric.next_control_state_0, non_ip_over_fabric_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, native_packet_over_fabric.next_control_state_1, ipv4_over_fabric_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, native_packet_over_fabric.next_control_state_2, ipv6_over_fabric_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, nexthop.next_control_state_0, nop_19.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, nexthop.next_control_state_1, set_nexthop_details_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, nexthop.next_control_state_2, set_nexthop_details_for_post_routed_flood_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv4_multicast.next_control_state_0, nop_20.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv4_multicast.next_control_state_1, on_miss_13.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv4_multicast.next_control_state_2, outer_multicast_route_s_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv4_multicast.next_control_state_3, outer_multicast_bridge_s_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv4_multicast_star_g.next_control_state_0, nop_21.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv4_multicast_star_g.next_control_state_1, outer_multicast_route_sm_star_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv4_multicast_star_g.next_control_state_2, outer_multicast_route_bidir_star_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv4_multicast_star_g.next_control_state_3, outer_multicast_bridge_star_g_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv6_multicast.next_control_state_0, nop_22.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv6_multicast.next_control_state_1, on_miss_14.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv6_multicast.next_control_state_2, outer_multicast_route_s_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv6_multicast.next_control_state_3, outer_multicast_bridge_s_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv6_multicast_star_g.next_control_state_0, nop_23.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv6_multicast_star_g.next_control_state_1, outer_multicast_route_sm_star_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv6_multicast_star_g.next_control_state_2, outer_multicast_route_bidir_star_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_ipv6_multicast_star_g.next_control_state_3, outer_multicast_bridge_star_g_hit_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_rmac.next_control_state_0, on_miss_15.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, outer_rmac.next_control_state_1, outer_rmac_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, port_vlan_mapping.next_control_state_0, set_bd_properties_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, port_vlan_mapping.next_control_state_1, port_vlan_mapping_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, qos.next_control_state_0, nop_24.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, qos.next_control_state_1, apply_cos_marking_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, qos.next_control_state_2, apply_dscp_marking_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, qos.next_control_state_3, apply_tc_marking_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rmac.next_control_state_0, rmac_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rmac.next_control_state_1, rmac_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, sflow_ing_take_sample.next_control_state_0, nop_25.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, sflow_ing_take_sample.next_control_state_1, sflow_ing_pkt_to_cpu_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, sflow_ingress.next_control_state_0, nop_26.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, sflow_ingress.next_control_state_1, sflow_ing_session_enable_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, smac.next_control_state_0, nop_27.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, smac.next_control_state_1, smac_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, smac.next_control_state_2, smac_hit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, spanning_tree.next_control_state_0, set_stp_state_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, storm_control.next_control_state_0, nop_28.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, storm_control.next_control_state_1, set_storm_control_meter_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, storm_control_stats.next_control_state_0, nop_29.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, switch_config_params.next_control_state_0, set_config_parameters_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, system_acl.next_control_state_0, nop_30.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, system_acl.next_control_state_1, redirect_to_cpu_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, system_acl.next_control_state_2, copy_to_cpu_with_reason_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, system_acl.next_control_state_3, copy_to_cpu_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, system_acl.next_control_state_4, drop_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, system_acl.next_control_state_5, drop_packet_with_reason_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, system_acl.next_control_state_6, negative_mirror_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel.next_control_state_0, nop_31.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel.next_control_state_1, tunnel_lookup_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel.next_control_state_2, terminate_tunnel_inner_non_ip_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel.next_control_state_3, terminate_tunnel_inner_ethernet_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel.next_control_state_4, terminate_tunnel_inner_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel.next_control_state_5, terminate_tunnel_inner_ethernet_ipv6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel.next_control_state_6, terminate_tunnel_inner_ipv6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_lookup_miss.next_control_state_0, non_ip_tunnel_lookup_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_lookup_miss.next_control_state_1, ipv4_tunnel_lookup_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_lookup_miss.next_control_state_2, ipv6_tunnel_lookup_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_miss.next_control_state_0, non_ip_tunnel_lookup_miss_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_miss.next_control_state_1, ipv4_tunnel_lookup_miss_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_miss.next_control_state_2, ipv6_tunnel_lookup_miss_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, urpf_bd.next_control_state_0, nop_32.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, urpf_bd.next_control_state_1, urpf_bd_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_mpls_packet.next_control_state_0, set_valid_mpls_label1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_mpls_packet.next_control_state_1, set_valid_mpls_label2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_mpls_packet.next_control_state_2, set_valid_mpls_label3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_0, malformed_outer_ethernet_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_1, set_valid_outer_unicast_packet_untagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_2, set_valid_outer_unicast_packet_single_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_3, set_valid_outer_unicast_packet_double_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_4, set_valid_outer_unicast_packet_qinq_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_5, set_valid_outer_multicast_packet_untagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_6, set_valid_outer_multicast_packet_single_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_7, set_valid_outer_multicast_packet_double_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_8, set_valid_outer_multicast_packet_qinq_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_9, set_valid_outer_broadcast_packet_untagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_10, set_valid_outer_broadcast_packet_single_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_11, set_valid_outer_broadcast_packet_double_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ethernet.next_control_state_12, set_valid_outer_broadcast_packet_qinq_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ipv4_packet.next_control_state_0, set_valid_outer_ipv4_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ipv4_packet.next_control_state_1, set_malformed_outer_ipv4_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ipv6_packet.next_control_state_0, set_valid_outer_ipv6_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_outer_ipv6_packet.next_control_state_1, set_malformed_outer_ipv6_packet_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_packet.next_control_state_0, nop_33.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_packet.next_control_state_1, set_unicast_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_packet.next_control_state_2, set_unicast_and_ipv6_src_is_link_local_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_packet.next_control_state_3, set_multicast_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_packet.next_control_state_4, set_multicast_and_ipv6_src_is_link_local_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_packet.next_control_state_5, set_broadcast_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, validate_packet.next_control_state_6, set_malformed_packet_0.prev_control_state);
  rule default_next_state if (default_req_ff.notEmpty);
    default_req_ff.deq;
    let _req = default_req_ff.first;
    let meta = _req.meta;
    let pkt = _req.pkt;
    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
    ingress_port_mapping_req_ff.enq(req);
  endrule

  rule acl_stats_next_state if (acl_stats_rsp_ff.notEmpty);
    acl_stats_rsp_ff.deq;
    let _rsp = acl_stats_rsp_ff.first;
    case (_rsp) matches
      tagged AclStatsAclStatsUpdateRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        storm_control_stats_req_ff.enq(req);
      end
    endcase
  endrule

  rule bd_flood_next_state if (bd_flood_rsp_ff.notEmpty);
    bd_flood_rsp_ff.deq;
    let _rsp = bd_flood_rsp_ff.first;
    case (_rsp) matches
      tagged BdFloodNopRspT {meta: .meta, pkt: .pkt}: begin
        let l2_metadata$learning_enabled = fromMaybe(?, meta.l2_metadata$learning_enabled);
        if (( l2_metadata$learning_enabled == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          learn_notify_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_lag_req_ff.enq(req);
        end
      end
      tagged BdFloodSetBdFloodMcIndexRspT {meta: .meta, pkt: .pkt}: begin
        let l2_metadata$learning_enabled = fromMaybe(?, meta.l2_metadata$learning_enabled);
        if (( l2_metadata$learning_enabled == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          learn_notify_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_lag_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule compute_ipv4_hashes_next_state if (compute_ipv4_hashes_rsp_ff.notEmpty);
    compute_ipv4_hashes_rsp_ff.deq;
    let _rsp = compute_ipv4_hashes_rsp_ff.first;
    case (_rsp) matches
      tagged ComputeIpv4HashesComputeLkpIpv4HashRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        compute_other_hashes_req_ff.enq(req);
      end
    endcase
  endrule

  rule compute_ipv6_hashes_next_state if (compute_ipv6_hashes_rsp_ff.notEmpty);
    compute_ipv6_hashes_rsp_ff.deq;
    let _rsp = compute_ipv6_hashes_rsp_ff.first;
    case (_rsp) matches
      tagged ComputeIpv6HashesComputeLkpIpv6HashRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        compute_other_hashes_req_ff.enq(req);
      end
    endcase
  endrule

  rule compute_non_ip_hashes_next_state if (compute_non_ip_hashes_rsp_ff.notEmpty);
    compute_non_ip_hashes_rsp_ff.deq;
    let _rsp = compute_non_ip_hashes_rsp_ff.first;
    case (_rsp) matches
      tagged ComputeNonIpHashesComputeLkpNonIpHashRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        compute_other_hashes_req_ff.enq(req);
      end
    endcase
  endrule

  rule compute_other_hashes_next_state if (compute_other_hashes_rsp_ff.notEmpty);
    compute_other_hashes_rsp_ff.deq;
    let _rsp = compute_other_hashes_rsp_ff.first;
    case (_rsp) matches
      tagged ComputeOtherHashesComputedTwoHashesRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_action_req_ff.enq(req);
        end
        else begin
          if (( ingress_metadata$port_type != 'h1 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            ingress_bd_stats_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            fabric_lag_req_ff.enq(req);
          end
        end
      end
      tagged ComputeOtherHashesComputedOneHashRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_action_req_ff.enq(req);
        end
        else begin
          if (( ingress_metadata$port_type != 'h1 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            ingress_bd_stats_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            fabric_lag_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule dmac_next_state if (dmac_rsp_ff.notEmpty);
    dmac_rsp_ff.deq;
    let _rsp = dmac_rsp_ff.first;
    case (_rsp) matches
      tagged DmacNopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        if (( l3_metadata$lkp_ip_type == 'h0 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            mac_acl_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            if (( l3_metadata$lkp_ip_type == 'h1 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ip_acl_req_ff.enq(req);
            end
            else begin
              if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ipv6_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
      end
      tagged DmacDmacHitRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        if (( l3_metadata$lkp_ip_type == 'h0 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            mac_acl_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            if (( l3_metadata$lkp_ip_type == 'h1 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ip_acl_req_ff.enq(req);
            end
            else begin
              if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ipv6_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
      end
      tagged DmacDmacMulticastHitRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        if (( l3_metadata$lkp_ip_type == 'h0 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            mac_acl_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            if (( l3_metadata$lkp_ip_type == 'h1 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ip_acl_req_ff.enq(req);
            end
            else begin
              if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ipv6_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
      end
      tagged DmacDmacMissRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        if (( l3_metadata$lkp_ip_type == 'h0 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            mac_acl_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            if (( l3_metadata$lkp_ip_type == 'h1 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ip_acl_req_ff.enq(req);
            end
            else begin
              if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ipv6_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
      end
      tagged DmacDmacRedirectNexthopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        if (( l3_metadata$lkp_ip_type == 'h0 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            mac_acl_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            if (( l3_metadata$lkp_ip_type == 'h1 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ip_acl_req_ff.enq(req);
            end
            else begin
              if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ipv6_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
      end
      tagged DmacDmacRedirectEcmpRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        if (( l3_metadata$lkp_ip_type == 'h0 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            mac_acl_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            if (( l3_metadata$lkp_ip_type == 'h1 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ip_acl_req_ff.enq(req);
            end
            else begin
              if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ipv6_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
      end
      tagged DmacDmacDropRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        if (( l3_metadata$lkp_ip_type == 'h0 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            mac_acl_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
            if (( l3_metadata$lkp_ip_type == 'h1 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ip_acl_req_ff.enq(req);
            end
            else begin
              if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ipv6_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            qos_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule drop_stats_next_state if (drop_stats_rsp_ff.notEmpty);
    drop_stats_rsp_ff.deq;
    let _rsp = drop_stats_rsp_ff.first;
    case (_rsp) matches
      tagged DropStatsDropStatsUpdateRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        next_req_ff.enq(req);
      end
    endcase
  endrule

  rule ecmp_group_next_state if (ecmp_group_rsp_ff.notEmpty);
    ecmp_group_rsp_ff.deq;
    let _rsp = ecmp_group_rsp_ff.first;
    case (_rsp) matches
      tagged EcmpGroupNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$egress_ifindex = fromMaybe(?, meta.ingress_metadata$egress_ifindex);
        if (( ingress_metadata$egress_ifindex == 'hffff )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          bd_flood_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          lag_group_req_ff.enq(req);
        end
      end
      tagged EcmpGroupSetEcmpNexthopDetailsRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$egress_ifindex = fromMaybe(?, meta.ingress_metadata$egress_ifindex);
        if (( ingress_metadata$egress_ifindex == 'hffff )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          bd_flood_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          lag_group_req_ff.enq(req);
        end
      end
      tagged EcmpGroupSetEcmpNexthopDetailsForPostRoutedFloodRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$egress_ifindex = fromMaybe(?, meta.ingress_metadata$egress_ifindex);
        if (( ingress_metadata$egress_ifindex == 'hffff )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          bd_flood_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          lag_group_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule fabric_ingress_dst_lkp_next_state if (fabric_ingress_dst_lkp_rsp_ff.notEmpty);
    fabric_ingress_dst_lkp_rsp_ff.deq;
    let _rsp = fabric_ingress_dst_lkp_rsp_ff.first;
    case (_rsp) matches
      tagged FabricIngressDstLkpNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type == 'h1 )) begin
          if (( isValid ( meta.valid_fabric_header_multicast ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            fabric_ingress_src_lkp_req_ff.enq(req);
          end
          else begin
            if (( tunnel_metadata$tunnel_terminate == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              native_packet_over_fabric_req_ff.enq(req);
            end
            else begin
              if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                outer_rmac_req_ff.enq(req);
              end
              else begin
                if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_miss_req_ff.enq(req);
                end
              end
            end
          end
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged FabricIngressDstLkpTerminateCpuPacketRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type == 'h1 )) begin
          if (( isValid ( meta.valid_fabric_header_multicast ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            fabric_ingress_src_lkp_req_ff.enq(req);
          end
          else begin
            if (( tunnel_metadata$tunnel_terminate == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              native_packet_over_fabric_req_ff.enq(req);
            end
            else begin
              if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                outer_rmac_req_ff.enq(req);
              end
              else begin
                if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_miss_req_ff.enq(req);
                end
              end
            end
          end
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged FabricIngressDstLkpSwitchFabricUnicastPacketRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type == 'h1 )) begin
          if (( isValid ( meta.valid_fabric_header_multicast ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            fabric_ingress_src_lkp_req_ff.enq(req);
          end
          else begin
            if (( tunnel_metadata$tunnel_terminate == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              native_packet_over_fabric_req_ff.enq(req);
            end
            else begin
              if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                outer_rmac_req_ff.enq(req);
              end
              else begin
                if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_miss_req_ff.enq(req);
                end
              end
            end
          end
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged FabricIngressDstLkpTerminateFabricUnicastPacketRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type == 'h1 )) begin
          if (( isValid ( meta.valid_fabric_header_multicast ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            fabric_ingress_src_lkp_req_ff.enq(req);
          end
          else begin
            if (( tunnel_metadata$tunnel_terminate == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              native_packet_over_fabric_req_ff.enq(req);
            end
            else begin
              if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                outer_rmac_req_ff.enq(req);
              end
              else begin
                if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_miss_req_ff.enq(req);
                end
              end
            end
          end
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged FabricIngressDstLkpSwitchFabricMulticastPacketRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type == 'h1 )) begin
          if (( isValid ( meta.valid_fabric_header_multicast ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            fabric_ingress_src_lkp_req_ff.enq(req);
          end
          else begin
            if (( tunnel_metadata$tunnel_terminate == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              native_packet_over_fabric_req_ff.enq(req);
            end
            else begin
              if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                outer_rmac_req_ff.enq(req);
              end
              else begin
                if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_miss_req_ff.enq(req);
                end
              end
            end
          end
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged FabricIngressDstLkpTerminateFabricMulticastPacketRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type == 'h1 )) begin
          if (( isValid ( meta.valid_fabric_header_multicast ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            fabric_ingress_src_lkp_req_ff.enq(req);
          end
          else begin
            if (( tunnel_metadata$tunnel_terminate == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              native_packet_over_fabric_req_ff.enq(req);
            end
            else begin
              if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                outer_rmac_req_ff.enq(req);
              end
              else begin
                if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  tunnel_miss_req_ff.enq(req);
                end
              end
            end
          end
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule fabric_ingress_src_lkp_next_state if (fabric_ingress_src_lkp_rsp_ff.notEmpty);
    fabric_ingress_src_lkp_rsp_ff.deq;
    let _rsp = fabric_ingress_src_lkp_rsp_ff.first;
    case (_rsp) matches
      tagged FabricIngressSrcLkpNopRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( tunnel_metadata$tunnel_terminate == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          native_packet_over_fabric_req_ff.enq(req);
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged FabricIngressSrcLkpSetIngressIfindexPropertiesRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( tunnel_metadata$tunnel_terminate == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          native_packet_over_fabric_req_ff.enq(req);
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule fabric_lag_next_state if (fabric_lag_rsp_ff.notEmpty);
    fabric_lag_rsp_ff.deq;
    let _rsp = fabric_lag_rsp_ff.first;
    case (_rsp) matches
      tagged FabricLagNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        if (( ingress_metadata$port_type != 'h1 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h20 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            system_acl_req_ff.enq(req);
          end
        end
      end
      tagged FabricLagSetFabricLagPortRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        if (( ingress_metadata$port_type != 'h1 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h20 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            system_acl_req_ff.enq(req);
          end
        end
      end
      tagged FabricLagSetFabricMulticastRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        if (( ingress_metadata$port_type != 'h1 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h20 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            system_acl_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule fwd_result_next_state if (fwd_result_rsp_ff.notEmpty);
    fwd_result_rsp_ff.deq;
    let _rsp = fwd_result_rsp_ff.first;
    case (_rsp) matches
      tagged FwdResultNopRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetL2RedirectActionRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetFibRedirectActionRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetCpuRedirectActionRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetAclRedirectActionRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetRaclRedirectActionRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetMulticastRouteActionRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetMulticastBridgeActionRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetMulticastFloodRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
      tagged FwdResultSetMulticastDropRspT {meta: .meta, pkt: .pkt}: begin
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( nexthop_metadata$nexthop_type == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ecmp_group_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          nexthop_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule ingress_bd_stats_next_state if (ingress_bd_stats_rsp_ff.notEmpty);
    ingress_bd_stats_rsp_ff.deq;
    let _rsp = ingress_bd_stats_rsp_ff.first;
    case (_rsp) matches
      tagged IngressBdStatsUpdateIngressBdStatsRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        acl_stats_req_ff.enq(req);
      end
    endcase
  endrule

  rule ingress_port_mapping_next_state if (ingress_port_mapping_rsp_ff.notEmpty);
    ingress_port_mapping_rsp_ff.deq;
    let _rsp = ingress_port_mapping_rsp_ff.first;
    case (_rsp) matches
      tagged IngressPortMappingSetIfindexRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ingress_port_properties_req_ff.enq(req);
      end
    endcase
  endrule

  rule ingress_port_properties_next_state if (ingress_port_properties_rsp_ff.notEmpty);
    ingress_port_properties_rsp_ff.deq;
    let _rsp = ingress_port_properties_rsp_ff.first;
    case (_rsp) matches
      tagged IngressPortPropertiesSetIngressPortPropertiesRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        validate_outer_ethernet_req_ff.enq(req);
      end
    endcase
  endrule

  rule int_sink_update_outer_next_state if (int_sink_update_outer_rsp_ff.notEmpty);
    int_sink_update_outer_rsp_ff.deq;
    let _rsp = int_sink_update_outer_rsp_ff.first;
    case (_rsp) matches
      tagged IntSinkUpdateOuterIntSinkUpdateVxlanGpeV4RspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_ingress_dst_lkp_req_ff.enq(req);
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged IntSinkUpdateOuterNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_ingress_dst_lkp_req_ff.enq(req);
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule int_source_next_state if (int_source_rsp_ff.notEmpty);
    int_source_rsp_ff.deq;
    let _rsp = int_source_rsp_ff.first;
    case (_rsp) matches
      tagged IntSourceIntSetSrcRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_ingress_dst_lkp_req_ff.enq(req);
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged IntSourceIntSetNoSrcRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( ingress_metadata$port_type != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_ingress_dst_lkp_req_ff.enq(req);
        end
        else begin
          if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_rmac_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule int_terminate_next_state if (int_terminate_rsp_ff.notEmpty);
    int_terminate_rsp_ff.deq;
    let _rsp = int_terminate_rsp_ff.first;
    case (_rsp) matches
      tagged IntTerminateIntSinkGpeRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_sink_update_outer_req_ff.enq(req);
      end
      tagged IntTerminateIntNoSinkRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_sink_update_outer_req_ff.enq(req);
      end
    endcase
  endrule

  rule ip_acl_next_state if (ip_acl_rsp_ff.notEmpty);
    ip_acl_rsp_ff.deq;
    let _rsp = ip_acl_rsp_ff.first;
    case (_rsp) matches
      tagged IpAclNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged IpAclAclDenyRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged IpAclAclPermitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged IpAclAclMirrorRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged IpAclAclRedirectNexthopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged IpAclAclRedirectEcmpRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
    endcase
  endrule

  rule ipsg_next_state if (ipsg_rsp_ff.notEmpty);
    ipsg_rsp_ff.deq;
    let _rsp = ipsg_rsp_ff.first;
    case (_rsp) matches
      tagged IpsgOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipsg_permit_special_req_ff.enq(req);
      end
    endcase
  endrule

  rule ipsg_permit_special_next_state if (ipsg_permit_special_rsp_ff.notEmpty);
    ipsg_permit_special_rsp_ff.deq;
    let _rsp = ipsg_permit_special_rsp_ff.first;
    case (_rsp) matches
      tagged IpsgPermitSpecialIpsgMissRspT {meta: .meta, pkt: .pkt}: begin
        if (( ! ( isValid ( meta.valid_int_header ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          int_source_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          int_terminate_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule ipv4_dest_vtep_next_state if (ipv4_dest_vtep_rsp_ff.notEmpty);
    ipv4_dest_vtep_rsp_ff.deq;
    let _rsp = ipv4_dest_vtep_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4DestVtepNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged Ipv4DestVtepSetTunnelTerminationFlagRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged Ipv4DestVtepSetTunnelVniAndTerminationFlagRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule ipv4_fib_next_state if (ipv4_fib_rsp_ff.notEmpty);
    ipv4_fib_rsp_ff.deq;
    let _rsp = ipv4_fib_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4FibOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv4_fib_lpm_req_ff.enq(req);
      end
      tagged Ipv4FibFibHitNexthopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged Ipv4FibFibHitEcmpRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule ipv4_fib_lpm_next_state if (ipv4_fib_lpm_rsp_ff.notEmpty);
    ipv4_fib_lpm_rsp_ff.deq;
    let _rsp = ipv4_fib_lpm_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4FibLpmOnMissRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged Ipv4FibLpmFibHitNexthopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged Ipv4FibLpmFibHitEcmpRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule ipv4_multicast_bridge_next_state if (ipv4_multicast_bridge_rsp_ff.notEmpty);
    ipv4_multicast_bridge_rsp_ff.deq;
    let _rsp = ipv4_multicast_bridge_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4MulticastBridgeOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv4_multicast_bridge_star_g_req_ff.enq(req);
      end
      tagged Ipv4MulticastBridgeMulticastBridgeSGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$ipv4_multicast_enabled = fromMaybe(?, meta.multicast_metadata$ipv4_multicast_enabled);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 ) && ( multicast_metadata$ipv4_multicast_enabled == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_multicast_route_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule ipv4_multicast_bridge_star_g_next_state if (ipv4_multicast_bridge_star_g_rsp_ff.notEmpty);
    ipv4_multicast_bridge_star_g_rsp_ff.deq;
    let _rsp = ipv4_multicast_bridge_star_g_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4MulticastBridgeStarGNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$ipv4_multicast_enabled = fromMaybe(?, meta.multicast_metadata$ipv4_multicast_enabled);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 ) && ( multicast_metadata$ipv4_multicast_enabled == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_multicast_route_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged Ipv4MulticastBridgeStarGMulticastBridgeStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$ipv4_multicast_enabled = fromMaybe(?, meta.multicast_metadata$ipv4_multicast_enabled);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 ) && ( multicast_metadata$ipv4_multicast_enabled == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_multicast_route_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule ipv4_multicast_route_next_state if (ipv4_multicast_route_rsp_ff.notEmpty);
    ipv4_multicast_route_rsp_ff.deq;
    let _rsp = ipv4_multicast_route_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4MulticastRouteOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv4_multicast_route_star_g_req_ff.enq(req);
      end
      tagged Ipv4MulticastRouteMulticastRouteSGHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule ipv4_multicast_route_star_g_next_state if (ipv4_multicast_route_star_g_rsp_ff.notEmpty);
    ipv4_multicast_route_star_g_rsp_ff.deq;
    let _rsp = ipv4_multicast_route_star_g_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4MulticastRouteStarGMulticastRouteStarGMissRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
      tagged Ipv4MulticastRouteStarGMulticastRouteSmStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
      tagged Ipv4MulticastRouteStarGMulticastRouteBidirStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule ipv4_racl_next_state if (ipv4_racl_rsp_ff.notEmpty);
    ipv4_racl_rsp_ff.deq;
    let _rsp = ipv4_racl_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4RaclNopRspT {meta: .meta, pkt: .pkt}: begin
        let ipv4_metadata$ipv4_urpf_mode = fromMaybe(?, meta.ipv4_metadata$ipv4_urpf_mode);
        if (( ipv4_metadata$ipv4_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_fib_req_ff.enq(req);
        end
      end
      tagged Ipv4RaclRaclDenyRspT {meta: .meta, pkt: .pkt}: begin
        let ipv4_metadata$ipv4_urpf_mode = fromMaybe(?, meta.ipv4_metadata$ipv4_urpf_mode);
        if (( ipv4_metadata$ipv4_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_fib_req_ff.enq(req);
        end
      end
      tagged Ipv4RaclRaclPermitRspT {meta: .meta, pkt: .pkt}: begin
        let ipv4_metadata$ipv4_urpf_mode = fromMaybe(?, meta.ipv4_metadata$ipv4_urpf_mode);
        if (( ipv4_metadata$ipv4_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_fib_req_ff.enq(req);
        end
      end
      tagged Ipv4RaclRaclRedirectNexthopRspT {meta: .meta, pkt: .pkt}: begin
        let ipv4_metadata$ipv4_urpf_mode = fromMaybe(?, meta.ipv4_metadata$ipv4_urpf_mode);
        if (( ipv4_metadata$ipv4_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_fib_req_ff.enq(req);
        end
      end
      tagged Ipv4RaclRaclRedirectEcmpRspT {meta: .meta, pkt: .pkt}: begin
        let ipv4_metadata$ipv4_urpf_mode = fromMaybe(?, meta.ipv4_metadata$ipv4_urpf_mode);
        if (( ipv4_metadata$ipv4_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_fib_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule ipv4_src_vtep_next_state if (ipv4_src_vtep_rsp_ff.notEmpty);
    ipv4_src_vtep_rsp_ff.deq;
    let _rsp = ipv4_src_vtep_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4SrcVtepOnMissRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged Ipv4SrcVtepSrcVtepHitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv4_dest_vtep_req_ff.enq(req);
      end
    endcase
  endrule

  rule ipv4_urpf_next_state if (ipv4_urpf_rsp_ff.notEmpty);
    ipv4_urpf_rsp_ff.deq;
    let _rsp = ipv4_urpf_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4UrpfOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv4_urpf_lpm_req_ff.enq(req);
      end
      tagged Ipv4UrpfIpv4UrpfHitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv4_fib_req_ff.enq(req);
      end
    endcase
  endrule

  rule ipv4_urpf_lpm_next_state if (ipv4_urpf_lpm_rsp_ff.notEmpty);
    ipv4_urpf_lpm_rsp_ff.deq;
    let _rsp = ipv4_urpf_lpm_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv4UrpfLpmIpv4UrpfHitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv4_fib_req_ff.enq(req);
      end
      tagged Ipv4UrpfLpmUrpfMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv4_fib_req_ff.enq(req);
      end
    endcase
  endrule

  rule ipv6_acl_next_state if (ipv6_acl_rsp_ff.notEmpty);
    ipv6_acl_rsp_ff.deq;
    let _rsp = ipv6_acl_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6AclNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged Ipv6AclAclDenyRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged Ipv6AclAclPermitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged Ipv6AclAclMirrorRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged Ipv6AclAclRedirectNexthopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged Ipv6AclAclRedirectEcmpRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
    endcase
  endrule

  rule ipv6_dest_vtep_next_state if (ipv6_dest_vtep_rsp_ff.notEmpty);
    ipv6_dest_vtep_rsp_ff.deq;
    let _rsp = ipv6_dest_vtep_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6DestVtepNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged Ipv6DestVtepSetTunnelTerminationFlagRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged Ipv6DestVtepSetTunnelVniAndTerminationFlagRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule ipv6_fib_next_state if (ipv6_fib_rsp_ff.notEmpty);
    ipv6_fib_rsp_ff.deq;
    let _rsp = ipv6_fib_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6FibOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv6_fib_lpm_req_ff.enq(req);
      end
      tagged Ipv6FibFibHitNexthopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged Ipv6FibFibHitEcmpRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule ipv6_fib_lpm_next_state if (ipv6_fib_lpm_rsp_ff.notEmpty);
    ipv6_fib_lpm_rsp_ff.deq;
    let _rsp = ipv6_fib_lpm_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6FibLpmOnMissRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged Ipv6FibLpmFibHitNexthopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged Ipv6FibLpmFibHitEcmpRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          urpf_bd_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule ipv6_multicast_bridge_next_state if (ipv6_multicast_bridge_rsp_ff.notEmpty);
    ipv6_multicast_bridge_rsp_ff.deq;
    let _rsp = ipv6_multicast_bridge_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6MulticastBridgeOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv6_multicast_bridge_star_g_req_ff.enq(req);
      end
      tagged Ipv6MulticastBridgeMulticastBridgeSGHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$ipv6_multicast_enabled = fromMaybe(?, meta.multicast_metadata$ipv6_multicast_enabled);
        if (( ( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 ) && ( multicast_metadata$ipv6_multicast_enabled == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_multicast_route_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule ipv6_multicast_bridge_star_g_next_state if (ipv6_multicast_bridge_star_g_rsp_ff.notEmpty);
    ipv6_multicast_bridge_star_g_rsp_ff.deq;
    let _rsp = ipv6_multicast_bridge_star_g_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6MulticastBridgeStarGNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$ipv6_multicast_enabled = fromMaybe(?, meta.multicast_metadata$ipv6_multicast_enabled);
        if (( ( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 ) && ( multicast_metadata$ipv6_multicast_enabled == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_multicast_route_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged Ipv6MulticastBridgeStarGMulticastBridgeStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$ipv6_multicast_enabled = fromMaybe(?, meta.multicast_metadata$ipv6_multicast_enabled);
        if (( ( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 ) && ( multicast_metadata$ipv6_multicast_enabled == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_multicast_route_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule ipv6_multicast_route_next_state if (ipv6_multicast_route_rsp_ff.notEmpty);
    ipv6_multicast_route_rsp_ff.deq;
    let _rsp = ipv6_multicast_route_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6MulticastRouteOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv6_multicast_route_star_g_req_ff.enq(req);
      end
      tagged Ipv6MulticastRouteMulticastRouteSGHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule ipv6_multicast_route_star_g_next_state if (ipv6_multicast_route_star_g_rsp_ff.notEmpty);
    ipv6_multicast_route_star_g_rsp_ff.deq;
    let _rsp = ipv6_multicast_route_star_g_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6MulticastRouteStarGMulticastRouteStarGMissRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
      tagged Ipv6MulticastRouteStarGMulticastRouteSmStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
      tagged Ipv6MulticastRouteStarGMulticastRouteBidirStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule ipv6_racl_next_state if (ipv6_racl_rsp_ff.notEmpty);
    ipv6_racl_rsp_ff.deq;
    let _rsp = ipv6_racl_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6RaclNopRspT {meta: .meta, pkt: .pkt}: begin
        let ipv6_metadata$ipv6_urpf_mode = fromMaybe(?, meta.ipv6_metadata$ipv6_urpf_mode);
        if (( ipv6_metadata$ipv6_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_fib_req_ff.enq(req);
        end
      end
      tagged Ipv6RaclRaclDenyRspT {meta: .meta, pkt: .pkt}: begin
        let ipv6_metadata$ipv6_urpf_mode = fromMaybe(?, meta.ipv6_metadata$ipv6_urpf_mode);
        if (( ipv6_metadata$ipv6_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_fib_req_ff.enq(req);
        end
      end
      tagged Ipv6RaclRaclPermitRspT {meta: .meta, pkt: .pkt}: begin
        let ipv6_metadata$ipv6_urpf_mode = fromMaybe(?, meta.ipv6_metadata$ipv6_urpf_mode);
        if (( ipv6_metadata$ipv6_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_fib_req_ff.enq(req);
        end
      end
      tagged Ipv6RaclRaclRedirectNexthopRspT {meta: .meta, pkt: .pkt}: begin
        let ipv6_metadata$ipv6_urpf_mode = fromMaybe(?, meta.ipv6_metadata$ipv6_urpf_mode);
        if (( ipv6_metadata$ipv6_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_fib_req_ff.enq(req);
        end
      end
      tagged Ipv6RaclRaclRedirectEcmpRspT {meta: .meta, pkt: .pkt}: begin
        let ipv6_metadata$ipv6_urpf_mode = fromMaybe(?, meta.ipv6_metadata$ipv6_urpf_mode);
        if (( ipv6_metadata$ipv6_urpf_mode != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_urpf_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv6_fib_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule ipv6_src_vtep_next_state if (ipv6_src_vtep_rsp_ff.notEmpty);
    ipv6_src_vtep_rsp_ff.deq;
    let _rsp = ipv6_src_vtep_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6SrcVtepOnMissRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged Ipv6SrcVtepSrcVtepHitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv6_dest_vtep_req_ff.enq(req);
      end
    endcase
  endrule

  rule ipv6_urpf_next_state if (ipv6_urpf_rsp_ff.notEmpty);
    ipv6_urpf_rsp_ff.deq;
    let _rsp = ipv6_urpf_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6UrpfOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv6_urpf_lpm_req_ff.enq(req);
      end
      tagged Ipv6UrpfIpv6UrpfHitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv6_fib_req_ff.enq(req);
      end
    endcase
  endrule

  rule ipv6_urpf_lpm_next_state if (ipv6_urpf_lpm_rsp_ff.notEmpty);
    ipv6_urpf_lpm_rsp_ff.deq;
    let _rsp = ipv6_urpf_lpm_rsp_ff.first;
    case (_rsp) matches
      tagged Ipv6UrpfLpmIpv6UrpfHitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv6_fib_req_ff.enq(req);
      end
      tagged Ipv6UrpfLpmUrpfMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        ipv6_fib_req_ff.enq(req);
      end
    endcase
  endrule

  rule lag_group_next_state if (lag_group_rsp_ff.notEmpty);
    lag_group_rsp_ff.deq;
    let _rsp = lag_group_rsp_ff.first;
    case (_rsp) matches
      tagged LagGroupSetLagMissRspT {meta: .meta, pkt: .pkt}: begin
        let l2_metadata$learning_enabled = fromMaybe(?, meta.l2_metadata$learning_enabled);
        if (( l2_metadata$learning_enabled == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          learn_notify_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_lag_req_ff.enq(req);
        end
      end
      tagged LagGroupSetLagPortRspT {meta: .meta, pkt: .pkt}: begin
        let l2_metadata$learning_enabled = fromMaybe(?, meta.l2_metadata$learning_enabled);
        if (( l2_metadata$learning_enabled == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          learn_notify_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_lag_req_ff.enq(req);
        end
      end
      tagged LagGroupSetLagRemotePortRspT {meta: .meta, pkt: .pkt}: begin
        let l2_metadata$learning_enabled = fromMaybe(?, meta.l2_metadata$learning_enabled);
        if (( l2_metadata$learning_enabled == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          learn_notify_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_lag_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule learn_notify_next_state if (learn_notify_rsp_ff.notEmpty);
    learn_notify_rsp_ff.deq;
    let _rsp = learn_notify_rsp_ff.first;
    case (_rsp) matches
      tagged LearnNotifyNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        fabric_lag_req_ff.enq(req);
      end
      tagged LearnNotifyGenerateLearnNotifyRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        fabric_lag_req_ff.enq(req);
      end
    endcase
  endrule

  rule mac_acl_next_state if (mac_acl_rsp_ff.notEmpty);
    mac_acl_rsp_ff.deq;
    let _rsp = mac_acl_rsp_ff.first;
    case (_rsp) matches
      tagged MacAclNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged MacAclAclDenyRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged MacAclAclPermitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged MacAclAclMirrorRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged MacAclAclRedirectNexthopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
      tagged MacAclAclRedirectEcmpRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        qos_req_ff.enq(req);
      end
    endcase
  endrule

  rule meter_action_next_state if (meter_action_rsp_ff.notEmpty);
    meter_action_rsp_ff.deq;
    let _rsp = meter_action_rsp_ff.first;
    case (_rsp) matches
      tagged MeterActionMeterPermitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        if (( ingress_metadata$port_type != 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ingress_bd_stats_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_lag_req_ff.enq(req);
        end
      end
      tagged MeterActionMeterDenyRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        if (( ingress_metadata$port_type != 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ingress_bd_stats_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fabric_lag_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule meter_index_next_state if (meter_index_rsp_ff.notEmpty);
    meter_index_rsp_ff.deq;
    let _rsp = meter_index_rsp_ff.first;
    case (_rsp) matches
      tagged MeterIndexNopRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          compute_ipv4_hashes_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv6_hashes_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_non_ip_hashes_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule mpls_next_state if (mpls_rsp_ff.notEmpty);
    mpls_rsp_ff.deq;
    let _rsp = mpls_rsp_ff.first;
    case (_rsp) matches
      tagged MplsTerminateEomplsRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged MplsTerminateVplsRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged MplsTerminateIpv4OverMplsRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged MplsTerminateIpv6OverMplsRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged MplsTerminatePwRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged MplsForwardMplsRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule native_packet_over_fabric_next_state if (native_packet_over_fabric_rsp_ff.notEmpty);
    native_packet_over_fabric_rsp_ff.deq;
    let _rsp = native_packet_over_fabric_rsp_ff.first;
    case (_rsp) matches
      tagged NativePacketOverFabricNonIpOverFabricRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          outer_rmac_req_ff.enq(req);
        end
        else begin
          if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_miss_req_ff.enq(req);
          end
        end
      end
      tagged NativePacketOverFabricIpv4OverFabricRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          outer_rmac_req_ff.enq(req);
        end
        else begin
          if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_miss_req_ff.enq(req);
          end
        end
      end
      tagged NativePacketOverFabricIpv6OverFabricRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( tunnel_metadata$ingress_tunnel_type != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          outer_rmac_req_ff.enq(req);
        end
        else begin
          if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_miss_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule nexthop_next_state if (nexthop_rsp_ff.notEmpty);
    nexthop_rsp_ff.deq;
    let _rsp = nexthop_rsp_ff.first;
    case (_rsp) matches
      tagged NexthopNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$egress_ifindex = fromMaybe(?, meta.ingress_metadata$egress_ifindex);
        if (( ingress_metadata$egress_ifindex == 'hffff )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          bd_flood_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          lag_group_req_ff.enq(req);
        end
      end
      tagged NexthopSetNexthopDetailsRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$egress_ifindex = fromMaybe(?, meta.ingress_metadata$egress_ifindex);
        if (( ingress_metadata$egress_ifindex == 'hffff )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          bd_flood_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          lag_group_req_ff.enq(req);
        end
      end
      tagged NexthopSetNexthopDetailsForPostRoutedFloodRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$egress_ifindex = fromMaybe(?, meta.ingress_metadata$egress_ifindex);
        if (( ingress_metadata$egress_ifindex == 'hffff )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          bd_flood_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          lag_group_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule outer_ipv4_multicast_next_state if (outer_ipv4_multicast_rsp_ff.notEmpty);
    outer_ipv4_multicast_rsp_ff.deq;
    let _rsp = outer_ipv4_multicast_rsp_ff.first;
    case (_rsp) matches
      tagged OuterIpv4MulticastNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv4MulticastOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        outer_ipv4_multicast_star_g_req_ff.enq(req);
      end
      tagged OuterIpv4MulticastOuterMulticastRouteSGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv4MulticastOuterMulticastBridgeSGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule outer_ipv4_multicast_star_g_next_state if (outer_ipv4_multicast_star_g_rsp_ff.notEmpty);
    outer_ipv4_multicast_star_g_rsp_ff.deq;
    let _rsp = outer_ipv4_multicast_star_g_rsp_ff.first;
    case (_rsp) matches
      tagged OuterIpv4MulticastStarGNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv4MulticastStarGOuterMulticastRouteSmStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv4MulticastStarGOuterMulticastRouteBidirStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv4MulticastStarGOuterMulticastBridgeStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule outer_ipv6_multicast_next_state if (outer_ipv6_multicast_rsp_ff.notEmpty);
    outer_ipv6_multicast_rsp_ff.deq;
    let _rsp = outer_ipv6_multicast_rsp_ff.first;
    case (_rsp) matches
      tagged OuterIpv6MulticastNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv6MulticastOnMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        outer_ipv6_multicast_star_g_req_ff.enq(req);
      end
      tagged OuterIpv6MulticastOuterMulticastRouteSGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv6MulticastOuterMulticastBridgeSGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule outer_ipv6_multicast_star_g_next_state if (outer_ipv6_multicast_star_g_rsp_ff.notEmpty);
    outer_ipv6_multicast_star_g_rsp_ff.deq;
    let _rsp = outer_ipv6_multicast_star_g_rsp_ff.first;
    case (_rsp) matches
      tagged OuterIpv6MulticastStarGNopRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv6MulticastStarGOuterMulticastRouteSmStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv6MulticastStarGOuterMulticastRouteBidirStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
      tagged OuterIpv6MulticastStarGOuterMulticastBridgeStarGHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_miss_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule outer_rmac_next_state if (outer_rmac_rsp_ff.notEmpty);
    outer_rmac_rsp_ff.deq;
    let _rsp = outer_rmac_rsp_ff.first;
    case (_rsp) matches
      tagged OuterRmacOnMissRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          outer_ipv4_multicast_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            outer_ipv6_multicast_req_ff.enq(req);
          end
          else begin
            if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_miss_req_ff.enq(req);
            end
          end
        end
      end
      tagged OuterRmacOuterRmacHitRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$mcast_rpf_group = fromMaybe(?, meta.multicast_metadata$mcast_rpf_group);
        let multicast_metadata$outer_mcast_route_hit = fromMaybe(?, meta.multicast_metadata$outer_mcast_route_hit);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$outer_mcast_mode = fromMaybe(?, meta.multicast_metadata$outer_mcast_mode);
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipv4_src_vtep_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            ipv6_src_vtep_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              mpls_req_ff.enq(req);
            end
            else begin
              if (( ( tunnel_metadata$tunnel_terminate == 'h1 ) || ( ( multicast_metadata$outer_mcast_route_hit == 'h1 ) && ( ( ( multicast_metadata$outer_mcast_mode == 'h1 ) && ( multicast_metadata$mcast_rpf_group == 'h0 ) ) || ( ( multicast_metadata$outer_mcast_mode == 'h2 ) && ( multicast_metadata$mcast_rpf_group != 'h0 ) ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                tunnel_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                tunnel_miss_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule port_vlan_mapping_next_state if (port_vlan_mapping_rsp_ff.notEmpty);
    port_vlan_mapping_rsp_ff.deq;
    let _rsp = port_vlan_mapping_rsp_ff.first;
    case (_rsp) matches
      tagged PortVlanMappingSetBdPropertiesRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l2_metadata$stp_group = fromMaybe(?, meta.l2_metadata$stp_group);
        let security_metadata$ipsg_enabled = fromMaybe(?, meta.security_metadata$ipsg_enabled);
        if (( ( ingress_metadata$port_type == 'h0 ) && ( l2_metadata$stp_group != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          spanning_tree_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$port_type == 'h0 ) && ( security_metadata$ipsg_enabled == 'h1 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            ipsg_req_ff.enq(req);
          end
          else begin
            if (( ! ( isValid ( meta.valid_int_header ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              int_source_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              int_terminate_req_ff.enq(req);
            end
          end
        end
      end
      tagged PortVlanMappingPortVlanMappingMissRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l2_metadata$stp_group = fromMaybe(?, meta.l2_metadata$stp_group);
        let security_metadata$ipsg_enabled = fromMaybe(?, meta.security_metadata$ipsg_enabled);
        if (( ( ingress_metadata$port_type == 'h0 ) && ( l2_metadata$stp_group != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          spanning_tree_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$port_type == 'h0 ) && ( security_metadata$ipsg_enabled == 'h1 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            ipsg_req_ff.enq(req);
          end
          else begin
            if (( ! ( isValid ( meta.valid_int_header ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              int_source_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              int_terminate_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule qos_next_state if (qos_rsp_ff.notEmpty);
    qos_rsp_ff.deq;
    let _rsp = qos_rsp_ff.first;
    case (_rsp) matches
      tagged QosNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        rmac_req_ff.enq(req);
      end
      tagged QosApplyCosMarkingRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        rmac_req_ff.enq(req);
      end
      tagged QosApplyDscpMarkingRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        rmac_req_ff.enq(req);
      end
      tagged QosApplyTcMarkingRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        rmac_req_ff.enq(req);
      end
    endcase
  endrule

  rule rmac_next_state if (rmac_rsp_ff.notEmpty);
    rmac_rsp_ff.deq;
    let _rsp = rmac_rsp_ff.first;
    case (_rsp) matches
      tagged RmacRmacHitRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ipv6_metadata$ipv6_unicast_enabled = fromMaybe(?, meta.ipv6_metadata$ipv6_unicast_enabled);
        let l3_metadata$urpf_mode = fromMaybe(?, meta.l3_metadata$urpf_mode);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let l3_metadata$urpf_hit = fromMaybe(?, meta.l3_metadata$urpf_hit);
        let ipv4_metadata$ipv4_unicast_enabled = fromMaybe(?, meta.ipv4_metadata$ipv4_unicast_enabled);
        if (( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 )) begin
          if (( ( l3_metadata$lkp_ip_type == 'h1 ) && ( ipv4_metadata$ipv4_unicast_enabled == 'h1 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            ipv4_racl_req_ff.enq(req);
          end
          else begin
            if (( ( l3_metadata$lkp_ip_type == 'h2 ) && ( ipv6_metadata$ipv6_unicast_enabled == 'h1 ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ipv6_racl_req_ff.enq(req);
            end
            else begin
              if (( ( l3_metadata$urpf_mode == 'h2 ) && ( l3_metadata$urpf_hit == 'h1 ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                urpf_bd_req_ff.enq(req);
              end
              else begin
                if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  meter_index_req_ff.enq(req);
                end
                else begin
                  if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    compute_ipv4_hashes_req_ff.enq(req);
                  end
                  else begin
                    if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      compute_ipv6_hashes_req_ff.enq(req);
                    end
                    else begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      compute_non_ip_hashes_req_ff.enq(req);
                    end
                  end
                end
              end
            end
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged RmacRmacMissRspT {meta: .meta, pkt: .pkt}: begin
        let multicast_metadata$ipv4_multicast_enabled = fromMaybe(?, meta.multicast_metadata$ipv4_multicast_enabled);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let multicast_metadata$ipv6_multicast_enabled = fromMaybe(?, meta.multicast_metadata$ipv6_multicast_enabled);
        if (( l3_metadata$lkp_ip_type == 'h1 )) begin
          if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            ipv4_multicast_bridge_req_ff.enq(req);
          end
          else begin
            if (( ( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 ) && ( multicast_metadata$ipv4_multicast_enabled == 'h1 ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ipv4_multicast_route_req_ff.enq(req);
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                meter_index_req_ff.enq(req);
              end
              else begin
                if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_ipv4_hashes_req_ff.enq(req);
                end
                else begin
                  if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    compute_ipv6_hashes_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    compute_non_ip_hashes_req_ff.enq(req);
                  end
                end
              end
            end
          end
        end
        else begin
          if (( l3_metadata$lkp_ip_type == 'h2 )) begin
            if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              ipv6_multicast_bridge_req_ff.enq(req);
            end
            else begin
              if (( ( ( ingress_metadata$bypass_lookups & 'h2 ) == 'h0 ) && ( multicast_metadata$ipv6_multicast_enabled == 'h1 ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ipv6_multicast_route_req_ff.enq(req);
              end
              else begin
                if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  meter_index_req_ff.enq(req);
                end
                else begin
                  if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    compute_ipv4_hashes_req_ff.enq(req);
                  end
                  else begin
                    if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      compute_ipv6_hashes_req_ff.enq(req);
                    end
                    else begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      compute_non_ip_hashes_req_ff.enq(req);
                    end
                  end
                end
              end
            end
          end
          else begin
            if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              meter_index_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv4_hashes_req_ff.enq(req);
              end
              else begin
                if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_ipv6_hashes_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_non_ip_hashes_req_ff.enq(req);
                end
              end
            end
          end
        end
      end
    endcase
  endrule

  rule sflow_ing_take_sample_next_state if (sflow_ing_take_sample_rsp_ff.notEmpty);
    sflow_ing_take_sample_rsp_ff.deq;
    let _rsp = sflow_ing_take_sample_rsp_ff.first;
    case (_rsp) matches
      tagged SflowIngTakeSampleNopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$fib_hit = fromMaybe(?, meta.l3_metadata$fib_hit);
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          storm_control_req_ff.enq(req);
        end
        else begin
          if (( ingress_metadata$port_type != 'h1 )) begin
            if (( ! ( ( isValid ( meta.valid_mpls[0] ) ) && ( l3_metadata$fib_hit == 'h1 ) ) )) begin
              if (( ingress_metadata$drop_flag == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                validate_packet_req_ff.enq(req);
              end
              else begin
                if (( ingress_metadata$port_type == 'h0 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  smac_req_ff.enq(req);
                end
                else begin
                  if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    dmac_req_ff.enq(req);
                  end
                  else begin
                    if (( l3_metadata$lkp_ip_type == 'h0 )) begin
                      if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                        mac_acl_req_ff.enq(req);
                      end
                      else begin
                        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                        qos_req_ff.enq(req);
                      end
                    end
                    else begin
                      if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                        if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                          ip_acl_req_ff.enq(req);
                        end
                        else begin
                          if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                            ipv6_acl_req_ff.enq(req);
                          end
                          else begin
                            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                            qos_req_ff.enq(req);
                          end
                        end
                      end
                      else begin
                        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                        qos_req_ff.enq(req);
                      end
                    end
                  end
                end
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                meter_index_req_ff.enq(req);
              end
              else begin
                if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_ipv4_hashes_req_ff.enq(req);
                end
                else begin
                  if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    compute_ipv6_hashes_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    compute_non_ip_hashes_req_ff.enq(req);
                  end
                end
              end
            end
          end
          else begin
            if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              meter_index_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv4_hashes_req_ff.enq(req);
              end
              else begin
                if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_ipv6_hashes_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_non_ip_hashes_req_ff.enq(req);
                end
              end
            end
          end
        end
      end
      tagged SflowIngTakeSampleSflowIngPktToCpuRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$fib_hit = fromMaybe(?, meta.l3_metadata$fib_hit);
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          storm_control_req_ff.enq(req);
        end
        else begin
          if (( ingress_metadata$port_type != 'h1 )) begin
            if (( ! ( ( isValid ( meta.valid_mpls[0] ) ) && ( l3_metadata$fib_hit == 'h1 ) ) )) begin
              if (( ingress_metadata$drop_flag == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                validate_packet_req_ff.enq(req);
              end
              else begin
                if (( ingress_metadata$port_type == 'h0 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  smac_req_ff.enq(req);
                end
                else begin
                  if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    dmac_req_ff.enq(req);
                  end
                  else begin
                    if (( l3_metadata$lkp_ip_type == 'h0 )) begin
                      if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                        mac_acl_req_ff.enq(req);
                      end
                      else begin
                        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                        qos_req_ff.enq(req);
                      end
                    end
                    else begin
                      if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                        if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                          ip_acl_req_ff.enq(req);
                        end
                        else begin
                          if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                            ipv6_acl_req_ff.enq(req);
                          end
                          else begin
                            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                            qos_req_ff.enq(req);
                          end
                        end
                      end
                      else begin
                        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                        qos_req_ff.enq(req);
                      end
                    end
                  end
                end
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                meter_index_req_ff.enq(req);
              end
              else begin
                if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_ipv4_hashes_req_ff.enq(req);
                end
                else begin
                  if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    compute_ipv6_hashes_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    compute_non_ip_hashes_req_ff.enq(req);
                  end
                end
              end
            end
          end
          else begin
            if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              meter_index_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv4_hashes_req_ff.enq(req);
              end
              else begin
                if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_ipv6_hashes_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_non_ip_hashes_req_ff.enq(req);
                end
              end
            end
          end
        end
      end
    endcase
  endrule

  rule sflow_ingress_next_state if (sflow_ingress_rsp_ff.notEmpty);
    sflow_ingress_rsp_ff.deq;
    let _rsp = sflow_ingress_rsp_ff.first;
    case (_rsp) matches
      tagged SflowIngressNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ing_take_sample_req_ff.enq(req);
      end
      tagged SflowIngressSflowIngSessionEnableRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ing_take_sample_req_ff.enq(req);
      end
    endcase
  endrule

  rule smac_next_state if (smac_rsp_ff.notEmpty);
    smac_rsp_ff.deq;
    let _rsp = smac_rsp_ff.first;
    case (_rsp) matches
      tagged SmacNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          dmac_req_ff.enq(req);
        end
        else begin
          if (( l3_metadata$lkp_ip_type == 'h0 )) begin
            if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              mac_acl_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              qos_req_ff.enq(req);
            end
          end
          else begin
            if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
              if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ip_acl_req_ff.enq(req);
              end
              else begin
                if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ipv6_acl_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  qos_req_ff.enq(req);
                end
              end
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              qos_req_ff.enq(req);
            end
          end
        end
      end
      tagged SmacSmacMissRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          dmac_req_ff.enq(req);
        end
        else begin
          if (( l3_metadata$lkp_ip_type == 'h0 )) begin
            if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              mac_acl_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              qos_req_ff.enq(req);
            end
          end
          else begin
            if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
              if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ip_acl_req_ff.enq(req);
              end
              else begin
                if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ipv6_acl_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  qos_req_ff.enq(req);
                end
              end
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              qos_req_ff.enq(req);
            end
          end
        end
      end
      tagged SmacSmacHitRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          dmac_req_ff.enq(req);
        end
        else begin
          if (( l3_metadata$lkp_ip_type == 'h0 )) begin
            if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              mac_acl_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              qos_req_ff.enq(req);
            end
          end
          else begin
            if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
              if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                ip_acl_req_ff.enq(req);
              end
              else begin
                if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ipv6_acl_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  qos_req_ff.enq(req);
                end
              end
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              qos_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule spanning_tree_next_state if (spanning_tree_rsp_ff.notEmpty);
    spanning_tree_rsp_ff.deq;
    let _rsp = spanning_tree_rsp_ff.first;
    case (_rsp) matches
      tagged SpanningTreeSetStpStateRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let security_metadata$ipsg_enabled = fromMaybe(?, meta.security_metadata$ipsg_enabled);
        if (( ( ingress_metadata$port_type == 'h0 ) && ( security_metadata$ipsg_enabled == 'h1 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          ipsg_req_ff.enq(req);
        end
        else begin
          if (( ! ( isValid ( meta.valid_int_header ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            int_source_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            int_terminate_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule storm_control_next_state if (storm_control_rsp_ff.notEmpty);
    storm_control_rsp_ff.deq;
    let _rsp = storm_control_rsp_ff.first;
    case (_rsp) matches
      tagged StormControlNopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$fib_hit = fromMaybe(?, meta.l3_metadata$fib_hit);
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ingress_metadata$port_type != 'h1 )) begin
          if (( ! ( ( isValid ( meta.valid_mpls[0] ) ) && ( l3_metadata$fib_hit == 'h1 ) ) )) begin
            if (( ingress_metadata$drop_flag == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_packet_req_ff.enq(req);
            end
            else begin
              if (( ingress_metadata$port_type == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                smac_req_ff.enq(req);
              end
              else begin
                if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  dmac_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h0 )) begin
                    if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      mac_acl_req_ff.enq(req);
                    end
                    else begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      qos_req_ff.enq(req);
                    end
                  end
                  else begin
                    if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                      if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                        ip_acl_req_ff.enq(req);
                      end
                      else begin
                        if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                          ipv6_acl_req_ff.enq(req);
                        end
                        else begin
                          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                          qos_req_ff.enq(req);
                        end
                      end
                    end
                    else begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      qos_req_ff.enq(req);
                    end
                  end
                end
              end
            end
          end
          else begin
            if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              meter_index_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv4_hashes_req_ff.enq(req);
              end
              else begin
                if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_ipv6_hashes_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_non_ip_hashes_req_ff.enq(req);
                end
              end
            end
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged StormControlSetStormControlMeterRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$fib_hit = fromMaybe(?, meta.l3_metadata$fib_hit);
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ingress_metadata$port_type != 'h1 )) begin
          if (( ! ( ( isValid ( meta.valid_mpls[0] ) ) && ( l3_metadata$fib_hit == 'h1 ) ) )) begin
            if (( ingress_metadata$drop_flag == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_packet_req_ff.enq(req);
            end
            else begin
              if (( ingress_metadata$port_type == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                smac_req_ff.enq(req);
              end
              else begin
                if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  dmac_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h0 )) begin
                    if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      mac_acl_req_ff.enq(req);
                    end
                    else begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      qos_req_ff.enq(req);
                    end
                  end
                  else begin
                    if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                      if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                        ip_acl_req_ff.enq(req);
                      end
                      else begin
                        if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                          ipv6_acl_req_ff.enq(req);
                        end
                        else begin
                          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                          qos_req_ff.enq(req);
                        end
                      end
                    end
                    else begin
                      MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                      qos_req_ff.enq(req);
                    end
                  end
                end
              end
            end
          end
          else begin
            if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              meter_index_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv4_hashes_req_ff.enq(req);
              end
              else begin
                if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_ipv6_hashes_req_ff.enq(req);
                end
                else begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  compute_non_ip_hashes_req_ff.enq(req);
                end
              end
            end
          end
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            meter_index_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv4_hashes_req_ff.enq(req);
            end
            else begin
              if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_ipv6_hashes_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                compute_non_ip_hashes_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  rule storm_control_stats_next_state if (storm_control_stats_rsp_ff.notEmpty);
    storm_control_stats_rsp_ff.deq;
    let _rsp = storm_control_stats_rsp_ff.first;
    case (_rsp) matches
      tagged StormControlStatsNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let nexthop_metadata$nexthop_type = fromMaybe(?, meta.nexthop_metadata$nexthop_type);
        if (( ! ( ingress_metadata$bypass_lookups == 'hffff ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          fwd_result_req_ff.enq(req);
        end
        else begin
          if (( nexthop_metadata$nexthop_type == 'h1 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            ecmp_group_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            nexthop_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule switch_config_params_next_state if (switch_config_params_rsp_ff.notEmpty);
    switch_config_params_rsp_ff.deq;
    let _rsp = switch_config_params_rsp_ff.first;
    case (_rsp) matches
      tagged SwitchConfigParamsSetConfigParametersRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        port_vlan_mapping_req_ff.enq(req);
      end
    endcase
  endrule

  rule system_acl_next_state if (system_acl_rsp_ff.notEmpty);
    system_acl_rsp_ff.deq;
    let _rsp = system_acl_rsp_ff.first;
    case (_rsp) matches
      tagged SystemAclNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        if (( ingress_metadata$drop_flag == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          drop_stats_req_ff.enq(req);
        end
      end
      tagged SystemAclRedirectToCpuRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        if (( ingress_metadata$drop_flag == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          drop_stats_req_ff.enq(req);
        end
      end
      tagged SystemAclCopyToCpuWithReasonRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        if (( ingress_metadata$drop_flag == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          drop_stats_req_ff.enq(req);
        end
      end
      tagged SystemAclCopyToCpuRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        if (( ingress_metadata$drop_flag == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          drop_stats_req_ff.enq(req);
        end
      end
      tagged SystemAclDropPacketRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        if (( ingress_metadata$drop_flag == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          drop_stats_req_ff.enq(req);
        end
      end
      tagged SystemAclDropPacketWithReasonRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        if (( ingress_metadata$drop_flag == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          drop_stats_req_ff.enq(req);
        end
      end
      tagged SystemAclNegativeMirrorRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$drop_flag = fromMaybe(?, meta.ingress_metadata$drop_flag);
        if (( ingress_metadata$drop_flag == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          drop_stats_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule tunnel_next_state if (tunnel_rsp_ff.notEmpty);
    tunnel_rsp_ff.deq;
    let _rsp = tunnel_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelTunnelLookupMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_lookup_miss_req_ff.enq(req);
      end
      tagged TunnelTerminateTunnelInnerNonIpRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelTerminateTunnelInnerEthernetIpv4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelTerminateTunnelInnerIpv4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelTerminateTunnelInnerEthernetIpv6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelTerminateTunnelInnerIpv6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_lookup_miss_next_state if (tunnel_lookup_miss_rsp_ff.notEmpty);
    tunnel_lookup_miss_rsp_ff.deq;
    let _rsp = tunnel_lookup_miss_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelLookupMissNonIpTunnelLookupMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelLookupMissIpv4TunnelLookupMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelLookupMissIpv6TunnelLookupMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_miss_next_state if (tunnel_miss_rsp_ff.notEmpty);
    tunnel_miss_rsp_ff.deq;
    let _rsp = tunnel_miss_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelMissNonIpTunnelLookupMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelMissIpv4TunnelLookupMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
      tagged TunnelMissIpv6TunnelLookupMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        sflow_ingress_req_ff.enq(req);
      end
    endcase
  endrule

  rule urpf_bd_next_state if (urpf_bd_rsp_ff.notEmpty);
    urpf_bd_rsp_ff.deq;
    let _rsp = urpf_bd_rsp_ff.first;
    case (_rsp) matches
      tagged UrpfBdNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
      tagged UrpfBdUrpfBdMissRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        if (( ( ingress_metadata$bypass_lookups & 'h10 ) == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          meter_index_req_ff.enq(req);
        end
        else begin
          if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv4 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv4 ) ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            compute_ipv4_hashes_req_ff.enq(req);
          end
          else begin
            if (( ( ( tunnel_metadata$tunnel_terminate == 'h0 ) && ( isValid ( meta.valid_ipv6 ) ) ) || ( ( tunnel_metadata$tunnel_terminate == 'h1 ) && ( isValid ( meta.valid_inner_ipv6 ) ) ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_ipv6_hashes_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              compute_non_ip_hashes_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule validate_mpls_packet_next_state if (validate_mpls_packet_rsp_ff.notEmpty);
    validate_mpls_packet_rsp_ff.deq;
    let _rsp = validate_mpls_packet_rsp_ff.first;
    case (_rsp) matches
      tagged ValidateMplsPacketSetValidMplsLabel1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        switch_config_params_req_ff.enq(req);
      end
      tagged ValidateMplsPacketSetValidMplsLabel2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        switch_config_params_req_ff.enq(req);
      end
      tagged ValidateMplsPacketSetValidMplsLabel3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        switch_config_params_req_ff.enq(req);
      end
    endcase
  endrule

  rule validate_outer_ethernet_next_state if (validate_outer_ethernet_rsp_ff.notEmpty);
    validate_outer_ethernet_rsp_ff.deq;
    let _rsp = validate_outer_ethernet_rsp_ff.first;
    case (_rsp) matches
      tagged ValidateOuterEthernetMalformedOuterEthernetPacketRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        switch_config_params_req_ff.enq(req);
      end
      tagged ValidateOuterEthernetSetValidOuterUnicastPacketUntaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterUnicastPacketSingleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterUnicastPacketDoubleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterUnicastPacketQinqTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterMulticastPacketUntaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterMulticastPacketSingleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterMulticastPacketDoubleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterMulticastPacketQinqTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterBroadcastPacketUntaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterBroadcastPacketSingleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterBroadcastPacketDoubleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
      tagged ValidateOuterEthernetSetValidOuterBroadcastPacketQinqTaggedRspT {meta: .meta, pkt: .pkt}: begin
        if (( isValid ( meta.valid_ipv4 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          validate_outer_ipv4_packet_req_ff.enq(req);
        end
        else begin
          if (( isValid ( meta.valid_ipv6 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            validate_outer_ipv6_packet_req_ff.enq(req);
          end
          else begin
            if (( isValid ( meta.valid_mpls[0] ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              validate_mpls_packet_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              switch_config_params_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule validate_outer_ipv4_packet_next_state if (validate_outer_ipv4_packet_rsp_ff.notEmpty);
    validate_outer_ipv4_packet_rsp_ff.deq;
    let _rsp = validate_outer_ipv4_packet_rsp_ff.first;
    case (_rsp) matches
      tagged ValidateOuterIpv4PacketSetValidOuterIpv4PacketRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        switch_config_params_req_ff.enq(req);
      end
      tagged ValidateOuterIpv4PacketSetMalformedOuterIpv4PacketRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        switch_config_params_req_ff.enq(req);
      end
    endcase
  endrule

  rule validate_outer_ipv6_packet_next_state if (validate_outer_ipv6_packet_rsp_ff.notEmpty);
    validate_outer_ipv6_packet_rsp_ff.deq;
    let _rsp = validate_outer_ipv6_packet_rsp_ff.first;
    case (_rsp) matches
      tagged ValidateOuterIpv6PacketSetValidOuterIpv6PacketRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        switch_config_params_req_ff.enq(req);
      end
      tagged ValidateOuterIpv6PacketSetMalformedOuterIpv6PacketRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        switch_config_params_req_ff.enq(req);
      end
    endcase
  endrule

  rule validate_packet_next_state if (validate_packet_rsp_ff.notEmpty);
    validate_packet_rsp_ff.deq;
    let _rsp = validate_packet_rsp_ff.first;
    case (_rsp) matches
      tagged ValidatePacketNopRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          smac_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            dmac_req_ff.enq(req);
          end
          else begin
            if (( l3_metadata$lkp_ip_type == 'h0 )) begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                mac_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ip_acl_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    ipv6_acl_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    qos_req_ff.enq(req);
                  end
                end
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged ValidatePacketSetUnicastRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          smac_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            dmac_req_ff.enq(req);
          end
          else begin
            if (( l3_metadata$lkp_ip_type == 'h0 )) begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                mac_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ip_acl_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    ipv6_acl_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    qos_req_ff.enq(req);
                  end
                end
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged ValidatePacketSetUnicastAndIpv6SrcIsLinkLocalRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          smac_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            dmac_req_ff.enq(req);
          end
          else begin
            if (( l3_metadata$lkp_ip_type == 'h0 )) begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                mac_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ip_acl_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    ipv6_acl_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    qos_req_ff.enq(req);
                  end
                end
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged ValidatePacketSetMulticastRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          smac_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            dmac_req_ff.enq(req);
          end
          else begin
            if (( l3_metadata$lkp_ip_type == 'h0 )) begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                mac_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ip_acl_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    ipv6_acl_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    qos_req_ff.enq(req);
                  end
                end
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged ValidatePacketSetMulticastAndIpv6SrcIsLinkLocalRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          smac_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            dmac_req_ff.enq(req);
          end
          else begin
            if (( l3_metadata$lkp_ip_type == 'h0 )) begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                mac_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ip_acl_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    ipv6_acl_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    qos_req_ff.enq(req);
                  end
                end
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged ValidatePacketSetBroadcastRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          smac_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            dmac_req_ff.enq(req);
          end
          else begin
            if (( l3_metadata$lkp_ip_type == 'h0 )) begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                mac_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ip_acl_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    ipv6_acl_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    qos_req_ff.enq(req);
                  end
                end
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
        end
      end
      tagged ValidatePacketSetMalformedPacketRspT {meta: .meta, pkt: .pkt}: begin
        let ingress_metadata$bypass_lookups = fromMaybe(?, meta.ingress_metadata$bypass_lookups);
        let ingress_metadata$port_type = fromMaybe(?, meta.ingress_metadata$port_type);
        let l3_metadata$lkp_ip_type = fromMaybe(?, meta.l3_metadata$lkp_ip_type);
        if (( ingress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          smac_req_ff.enq(req);
        end
        else begin
          if (( ( ingress_metadata$bypass_lookups & 'h1 ) == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            dmac_req_ff.enq(req);
          end
          else begin
            if (( l3_metadata$lkp_ip_type == 'h0 )) begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                mac_acl_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
            else begin
              if (( ( ingress_metadata$bypass_lookups & 'h4 ) == 'h0 )) begin
                if (( l3_metadata$lkp_ip_type == 'h1 )) begin
                  MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                  ip_acl_req_ff.enq(req);
                end
                else begin
                  if (( l3_metadata$lkp_ip_type == 'h2 )) begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    ipv6_acl_req_ff.enq(req);
                  end
                  else begin
                    MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                    qos_req_ff.enq(req);
                  end
                end
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                qos_req_ff.enq(req);
              end
            end
          end
        end
      end
    endcase
  endrule

  interface next = (interface Client#(MetadataRequest, MetadataResponse);
    interface request = toGet(next_req_ff);
    interface response = toPut(next_rsp_ff);
  endinterface);
endmodule

// ====== EGRESS_ACL ======

typedef struct {
  Bit#(1) padding;
  Bit#(9) standard_metadata$egress_port;
  Bit#(1) intrinsic_metadata$deflection_flag;
  Bit#(16) l3_metadata$l3_mtu_check;
} EgressAclReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_EGRESS_ACL,
  NOP,
  EGRESS_MIRROR,
  EGRESS_MIRROR_DROP,
  EGRESS_REDIRECT_TO_CPU
} EgressAclActionT deriving (Bits, Eq, FShow);
typedef struct {
  EgressAclActionT _action;
  Bit#(32) runtime_session_id;
  Bit#(16) runtime_reason_code;
} EgressAclRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(51)) matchtable_read_egress_acl(Bit#(27) msgtype);
import "BDPI" function Action matchtable_write_egress_acl(Bit#(27) msgtype, Bit#(51) data);
`endif
instance MatchTableSim#(97, 27, 51);
  function ActionValue#(Bit#(51)) matchtable_read(Bit#(97) id, Bit#(27) key);
    actionvalue
      let v <- matchtable_read_egress_acl(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(97) id, Bit#(27) key, Bit#(51) data);
    action
      matchtable_write_egress_acl(key, data);
    endaction
  endfunction

endinstance
interface EgressAcl;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
endinterface
(* synthesize *)
module mkEgressAcl  (EgressAcl);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(4, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(4, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(97, 512, SizeOf#(EgressAclReqT), SizeOf#(EgressAclRspT)) matchTable <- mkMatchTable("egress_acl.dat");
  Vector#(4, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(4) readyChannel = -1;
  for (Integer i=3; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let standard_metadata$egress_port = fromMaybe(?, meta.standard_metadata$egress_port);
    let intrinsic_metadata$deflection_flag = fromMaybe(?, meta.intrinsic_metadata$deflection_flag);
    let l3_metadata$l3_mtu_check = fromMaybe(?, meta.l3_metadata$l3_mtu_check);
    EgressAclReqT req = EgressAclReqT {standard_metadata$egress_port: standard_metadata$egress_port,intrinsic_metadata$deflection_flag: intrinsic_metadata$deflection_flag,l3_metadata$l3_mtu_check: l3_metadata$l3_mtu_check};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      EgressAclRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        EGRESS_MIRROR: begin
          BBRequest req = tagged EgressMirrorReqT {pkt: pkt, runtime_session_id: resp.runtime_session_id};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        EGRESS_MIRROR_DROP: begin
          BBRequest req = tagged EgressMirrorDropReqT {pkt: pkt, runtime_session_id: resp.runtime_session_id};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        EGRESS_REDIRECT_TO_CPU: begin
          BBRequest req = tagged EgressRedirectToCpuReqT {pkt: pkt, runtime_reason_code: resp.runtime_reason_code};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged EgressAclNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged EgressMirrorRspT {pkt: .pkt, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id}: begin
        meta.i2e_metadata$mirror_session_id = tagged Valid i2e_metadata$mirror_session_id;
        MetadataResponse rsp = tagged EgressAclEgressMirrorRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged EgressMirrorDropRspT {pkt: .pkt, i2e_metadata$mirror_session_id: .i2e_metadata$mirror_session_id}: begin
        meta.i2e_metadata$mirror_session_id = tagged Valid i2e_metadata$mirror_session_id;
        MetadataResponse rsp = tagged EgressAclEgressMirrorDropRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged EgressRedirectToCpuRspT {pkt: .pkt, fabric_metadata$reason_code: .fabric_metadata$reason_code}: begin
        meta.fabric_metadata$reason_code = tagged Valid fabric_metadata$reason_code;
        MetadataResponse rsp = tagged EgressAclEgressRedirectToCpuRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
endmodule

// ====== EGRESS_BD_MAP ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) egress_metadata$bd;
} EgressBdMapReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_EGRESS_BD_MAP,
  NOP,
  SET_EGRESS_BD_PROPERTIES
} EgressBdMapActionT deriving (Bits, Eq, FShow);
typedef struct {
  EgressBdMapActionT _action;
  Bit#(9) runtime_smac_idx;
} EgressBdMapRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(11)) matchtable_read_egress_bd_map(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_egress_bd_map(Bit#(18) msgtype, Bit#(11) data);
`endif
instance MatchTableSim#(81, 18, 11);
  function ActionValue#(Bit#(11)) matchtable_read(Bit#(81) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_egress_bd_map(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(81) id, Bit#(18) key, Bit#(11) data);
    action
      matchtable_write_egress_bd_map(key, data);
    endaction
  endfunction

endinstance
interface EgressBdMap;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkEgressBdMap  (EgressBdMap);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(81, 1024, SizeOf#(EgressBdMapReqT), SizeOf#(EgressBdMapRspT)) matchTable <- mkMatchTable("egress_bd_map.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let egress_metadata$bd = fromMaybe(?, meta.egress_metadata$bd);
    EgressBdMapReqT req = EgressBdMapReqT {egress_metadata$bd: egress_metadata$bd};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      EgressBdMapRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_EGRESS_BD_PROPERTIES: begin
          BBRequest req = tagged SetEgressBdPropertiesReqT {pkt: pkt, runtime_smac_idx: resp.runtime_smac_idx};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged EgressBdMapNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetEgressBdPropertiesRspT {pkt: .pkt, egress_metadata$smac_idx: .egress_metadata$smac_idx}: begin
        meta.egress_metadata$smac_idx = tagged Valid egress_metadata$smac_idx;
        MetadataResponse rsp = tagged EgressBdMapSetEgressBdPropertiesRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== EGRESS_BD_STATS ======

typedef struct {
  Bit#(8) padding;
  Bit#(16) egress_metadata$bd;
  Bit#(3) l2_metadata$lkp_pkt_type;
} EgressBdStatsReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_EGRESS_BD_STATS,
  NOP
} EgressBdStatsActionT deriving (Bits, Eq, FShow);
typedef struct {
  EgressBdStatsActionT _action;
} EgressBdStatsRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_egress_bd_stats(Bit#(27) msgtype);
import "BDPI" function Action matchtable_write_egress_bd_stats(Bit#(27) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(80, 27, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(80) id, Bit#(27) key);
    actionvalue
      let v <- matchtable_read_egress_bd_stats(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(80) id, Bit#(27) key, Bit#(1) data);
    action
      matchtable_write_egress_bd_stats(key, data);
    endaction
  endfunction

endinstance
interface EgressBdStats;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkEgressBdStats  (EgressBdStats);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(80, 1024, SizeOf#(EgressBdStatsReqT), SizeOf#(EgressBdStatsRspT)) matchTable <- mkMatchTable("egress_bd_stats.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let egress_metadata$bd = fromMaybe(?, meta.egress_metadata$bd);
    let l2_metadata$lkp_pkt_type = fromMaybe(?, meta.l2_metadata$lkp_pkt_type);
    EgressBdStatsReqT req = EgressBdStatsReqT {egress_metadata$bd: egress_metadata$bd,l2_metadata$lkp_pkt_type: l2_metadata$lkp_pkt_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      EgressBdStatsRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged EgressBdStatsNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== EGRESS_FILTER ======

typedef struct {
} EgressFilterReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_EGRESS_FILTER,
  EGRESS_FILTER_CHECK
} EgressFilterActionT deriving (Bits, Eq, FShow);
typedef struct {
  EgressFilterActionT _action;
} EgressFilterRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_egress_filter(Bit#(0) msgtype);
import "BDPI" function Action matchtable_write_egress_filter(Bit#(0) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(103, 0, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(103) id, Bit#(0) key);
    actionvalue
      let v <- matchtable_read_egress_filter(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(103) id, Bit#(0) key, Bit#(1) data);
    action
      matchtable_write_egress_filter(key, data);
    endaction
  endfunction

endinstance
interface EgressFilter;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkEgressFilter  (EgressFilter);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  FIFOF#(MetadataT) metadata_ff <- mkFIFOF;
  rule rl_handle_action_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    packet_ff.enq(pkt);
    metadata_ff.enq(meta);
    BBRequest req = tagged EgressFilterCheckReqT {pkt: pkt};
    bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
  endrule

  rule rl_handle_action_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff).get;
    case (v) matches
      tagged EgressFilterCheckRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged EgressFilterEgressFilterCheckRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== EGRESS_FILTER_DROP ======

typedef struct {
} EgressFilterDropReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_EGRESS_FILTER_DROP,
  SET_EGRESS_FILTER_DROP
} EgressFilterDropActionT deriving (Bits, Eq, FShow);
typedef struct {
  EgressFilterDropActionT _action;
} EgressFilterDropRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_egress_filter_drop(Bit#(0) msgtype);
import "BDPI" function Action matchtable_write_egress_filter_drop(Bit#(0) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(102, 0, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(102) id, Bit#(0) key);
    actionvalue
      let v <- matchtable_read_egress_filter_drop(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(102) id, Bit#(0) key, Bit#(1) data);
    action
      matchtable_write_egress_filter_drop(key, data);
    endaction
  endfunction

endinstance
interface EgressFilterDrop;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkEgressFilterDrop  (EgressFilterDrop);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  FIFOF#(MetadataT) metadata_ff <- mkFIFOF;
  rule rl_handle_action_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    packet_ff.enq(pkt);
    metadata_ff.enq(meta);
    BBRequest req = tagged SetEgressFilterDropReqT {pkt: pkt};
    bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
  endrule

  rule rl_handle_action_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff).get;
    case (v) matches
      tagged SetEgressFilterDropRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged EgressFilterDropSetEgressFilterDropRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== EGRESS_PORT_MAPPING ======

typedef struct {
  Bit#(9) standard_metadata$egress_port;
} EgressPortMappingReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_EGRESS_PORT_MAPPING,
  EGRESS_PORT_TYPE_NORMAL,
  EGRESS_PORT_TYPE_FABRIC,
  EGRESS_PORT_TYPE_CPU
} EgressPortMappingActionT deriving (Bits, Eq, FShow);
typedef struct {
  EgressPortMappingActionT _action;
  Bit#(16) runtime_ifindex;
} EgressPortMappingRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_egress_port_mapping(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_egress_port_mapping(Bit#(9) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(78, 9, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(78) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_egress_port_mapping(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(78) id, Bit#(9) key, Bit#(18) data);
    action
      matchtable_write_egress_port_mapping(key, data);
    endaction
  endfunction

endinstance
interface EgressPortMapping;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkEgressPortMapping  (EgressPortMapping);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(78, 512, SizeOf#(EgressPortMappingReqT), SizeOf#(EgressPortMappingRspT)) matchTable <- mkMatchTable("egress_port_mapping.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let standard_metadata$egress_port = fromMaybe(?, meta.standard_metadata$egress_port);
    EgressPortMappingReqT req = EgressPortMappingReqT {standard_metadata$egress_port: standard_metadata$egress_port};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      EgressPortMappingRspT resp = unpack(data);
      case (resp._action) matches
        EGRESS_PORT_TYPE_NORMAL: begin
          BBRequest req = tagged EgressPortTypeNormalReqT {pkt: pkt, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        EGRESS_PORT_TYPE_FABRIC: begin
          BBRequest req = tagged EgressPortTypeFabricReqT {pkt: pkt, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        EGRESS_PORT_TYPE_CPU: begin
          BBRequest req = tagged EgressPortTypeCpuReqT {pkt: pkt, runtime_ifindex: resp.runtime_ifindex};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged EgressPortTypeNormalRspT {pkt: .pkt, egress_metadata$ifindex: .egress_metadata$ifindex, egress_metadata$port_type: .egress_metadata$port_type}: begin
        meta.egress_metadata$ifindex = tagged Valid egress_metadata$ifindex;
        meta.egress_metadata$port_type = tagged Valid egress_metadata$port_type;
        MetadataResponse rsp = tagged EgressPortMappingEgressPortTypeNormalRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged EgressPortTypeFabricRspT {pkt: .pkt, egress_metadata$ifindex: .egress_metadata$ifindex, egress_metadata$port_type: .egress_metadata$port_type, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type}: begin
        meta.egress_metadata$ifindex = tagged Valid egress_metadata$ifindex;
        meta.egress_metadata$port_type = tagged Valid egress_metadata$port_type;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        MetadataResponse rsp = tagged EgressPortMappingEgressPortTypeFabricRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged EgressPortTypeCpuRspT {pkt: .pkt, egress_metadata$ifindex: .egress_metadata$ifindex, egress_metadata$port_type: .egress_metadata$port_type, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type}: begin
        meta.egress_metadata$ifindex = tagged Valid egress_metadata$ifindex;
        meta.egress_metadata$port_type = tagged Valid egress_metadata$port_type;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        MetadataResponse rsp = tagged EgressPortMappingEgressPortTypeCpuRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== EGRESS_VLAN_XLATE ======

typedef struct {
  Bit#(4) padding;
  Bit#(16) egress_metadata$ifindex;
  Bit#(16) egress_metadata$bd;
} EgressVlanXlateReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_EGRESS_VLAN_XLATE,
  SET_EGRESS_PACKET_VLAN_UNTAGGED,
  SET_EGRESS_PACKET_VLAN_TAGGED,
  SET_EGRESS_PACKET_VLAN_DOUBLE_TAGGED
} EgressVlanXlateActionT deriving (Bits, Eq, FShow);
typedef struct {
  EgressVlanXlateActionT _action;
  Bit#(12) runtime_vlan_id;
  Bit#(12) runtime_s_tag;
  Bit#(12) runtime_c_tag;
} EgressVlanXlateRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(38)) matchtable_read_egress_vlan_xlate(Bit#(36) msgtype);
import "BDPI" function Action matchtable_write_egress_vlan_xlate(Bit#(36) msgtype, Bit#(38) data);
`endif
instance MatchTableSim#(79, 36, 38);
  function ActionValue#(Bit#(38)) matchtable_read(Bit#(79) id, Bit#(36) key);
    actionvalue
      let v <- matchtable_read_egress_vlan_xlate(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(79) id, Bit#(36) key, Bit#(38) data);
    action
      matchtable_write_egress_vlan_xlate(key, data);
    endaction
  endfunction

endinstance
interface EgressVlanXlate;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkEgressVlanXlate  (EgressVlanXlate);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(79, 1024, SizeOf#(EgressVlanXlateReqT), SizeOf#(EgressVlanXlateRspT)) matchTable <- mkMatchTable("egress_vlan_xlate.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let egress_metadata$ifindex = fromMaybe(?, meta.egress_metadata$ifindex);
    let egress_metadata$bd = fromMaybe(?, meta.egress_metadata$bd);
    EgressVlanXlateReqT req = EgressVlanXlateReqT {egress_metadata$ifindex: egress_metadata$ifindex,egress_metadata$bd: egress_metadata$bd};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      EgressVlanXlateRspT resp = unpack(data);
      case (resp._action) matches
        SET_EGRESS_PACKET_VLAN_UNTAGGED: begin
          BBRequest req = tagged SetEgressPacketVlanUntaggedReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_EGRESS_PACKET_VLAN_TAGGED: begin
          BBRequest req = tagged SetEgressPacketVlanTaggedReqT {pkt: pkt, ethernet$etherType: ethernet$etherType, runtime_vlan_id: resp.runtime_vlan_id};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_EGRESS_PACKET_VLAN_DOUBLE_TAGGED: begin
          BBRequest req = tagged SetEgressPacketVlanDoubleTaggedReqT {pkt: pkt, ethernet$etherType: ethernet$etherType, runtime_c_tag: resp.runtime_c_tag, runtime_s_tag: resp.runtime_s_tag};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged SetEgressPacketVlanUntaggedRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged EgressVlanXlateSetEgressPacketVlanUntaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetEgressPacketVlanTaggedRspT {pkt: .pkt, vlan_tag_0$vid: .vlan_tag_0$vid, vlan_tag_0$etherType: .vlan_tag_0$etherType, ethernet$etherType: .ethernet$etherType}: begin
        meta.vlan_tag_0$vid = tagged Valid vlan_tag_0$vid;
        meta.vlan_tag_0$etherType = tagged Valid vlan_tag_0$etherType;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged EgressVlanXlateSetEgressPacketVlanTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetEgressPacketVlanDoubleTaggedRspT {pkt: .pkt, vlan_tag_1$vid: .vlan_tag_1$vid, vlan_tag_0$vid: .vlan_tag_0$vid, vlan_tag_0$etherType: .vlan_tag_0$etherType, vlan_tag_1$etherType: .vlan_tag_1$etherType, ethernet$etherType: .ethernet$etherType}: begin
        meta.vlan_tag_1$vid = tagged Valid vlan_tag_1$vid;
        meta.vlan_tag_0$vid = tagged Valid vlan_tag_0$vid;
        meta.vlan_tag_0$etherType = tagged Valid vlan_tag_0$etherType;
        meta.vlan_tag_1$etherType = tagged Valid vlan_tag_1$etherType;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged EgressVlanXlateSetEgressPacketVlanDoubleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== EGRESS_VNI ======

typedef struct {
  Bit#(6) padding;
  Bit#(16) egress_metadata$bd;
  Bit#(5) tunnel_metadata$egress_tunnel_type;
} EgressVniReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_EGRESS_VNI,
  NOP,
  SET_EGRESS_TUNNEL_VNI
} EgressVniActionT deriving (Bits, Eq, FShow);
typedef struct {
  EgressVniActionT _action;
  Bit#(24) runtime_vnid;
} EgressVniRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(26)) matchtable_read_egress_vni(Bit#(27) msgtype);
import "BDPI" function Action matchtable_write_egress_vni(Bit#(27) msgtype, Bit#(26) data);
`endif
instance MatchTableSim#(88, 27, 26);
  function ActionValue#(Bit#(26)) matchtable_read(Bit#(88) id, Bit#(27) key);
    actionvalue
      let v <- matchtable_read_egress_vni(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(88) id, Bit#(27) key, Bit#(26) data);
    action
      matchtable_write_egress_vni(key, data);
    endaction
  endfunction

endinstance
interface EgressVni;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkEgressVni  (EgressVni);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(88, 1024, SizeOf#(EgressVniReqT), SizeOf#(EgressVniRspT)) matchTable <- mkMatchTable("egress_vni.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let egress_metadata$bd = fromMaybe(?, meta.egress_metadata$bd);
    let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
    EgressVniReqT req = EgressVniReqT {egress_metadata$bd: egress_metadata$bd,tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      EgressVniRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_EGRESS_TUNNEL_VNI: begin
          BBRequest req = tagged SetEgressTunnelVniReqT {pkt: pkt, runtime_vnid: resp.runtime_vnid};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged EgressVniNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetEgressTunnelVniRspT {pkt: .pkt, tunnel_metadata$vnid: .tunnel_metadata$vnid}: begin
        meta.tunnel_metadata$vnid = tagged Valid tunnel_metadata$vnid;
        MetadataResponse rsp = tagged EgressVniSetEgressTunnelVniRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== INT_BOS ======

typedef struct {
  Bit#(3) padding;
  Bit#(8) int_header$total_hop_cnt;
  Bit#(4) int_header$instruction_mask_0003;
  Bit#(4) int_header$instruction_mask_0407;
  Bit#(4) int_header$instruction_mask_0811;
  Bit#(4) int_header$instruction_mask_1215;
} IntBosReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_BOS,
  INT_SET_HEADER_0_BOS,
  INT_SET_HEADER_1_BOS,
  INT_SET_HEADER_2_BOS,
  INT_SET_HEADER_3_BOS,
  INT_SET_HEADER_4_BOS,
  INT_SET_HEADER_5_BOS,
  INT_SET_HEADER_6_BOS,
  INT_SET_HEADER_7_BOS,
  NOP
} IntBosActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntBosActionT _action;
} IntBosRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(4)) matchtable_read_int_bos(Bit#(27) msgtype);
import "BDPI" function Action matchtable_write_int_bos(Bit#(27) msgtype, Bit#(4) data);
`endif
instance MatchTableSim#(109, 27, 4);
  function ActionValue#(Bit#(4)) matchtable_read(Bit#(109) id, Bit#(27) key);
    actionvalue
      let v <- matchtable_read_int_bos(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(109) id, Bit#(27) key, Bit#(4) data);
    action
      matchtable_write_int_bos(key, data);
    endaction
  endfunction

endinstance
interface IntBos;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
endinterface
(* synthesize *)
module mkIntBos  (IntBos);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(9, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(9, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(109, 256, SizeOf#(IntBosReqT), SizeOf#(IntBosRspT)) matchTable <- mkMatchTable("int_bos.dat");
  Vector#(9, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(9) readyChannel = -1;
  for (Integer i=8; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let int_header$total_hop_cnt = fromMaybe(?, meta.int_header$total_hop_cnt);
    let int_header$instruction_mask_0003 = fromMaybe(?, meta.int_header$instruction_mask_0003);
    let int_header$instruction_mask_0407 = fromMaybe(?, meta.int_header$instruction_mask_0407);
    let int_header$instruction_mask_0811 = fromMaybe(?, meta.int_header$instruction_mask_0811);
    let int_header$instruction_mask_1215 = fromMaybe(?, meta.int_header$instruction_mask_1215);
    IntBosReqT req = IntBosReqT {int_header$total_hop_cnt: int_header$total_hop_cnt,int_header$instruction_mask_0003: int_header$instruction_mask_0003,int_header$instruction_mask_0407: int_header$instruction_mask_0407,int_header$instruction_mask_0811: int_header$instruction_mask_0811,int_header$instruction_mask_1215: int_header$instruction_mask_1215};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntBosRspT resp = unpack(data);
      case (resp._action) matches
        INT_SET_HEADER_0_BOS: begin
          BBRequest req = tagged IntSetHeader0BosReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_1_BOS: begin
          BBRequest req = tagged IntSetHeader1BosReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_2_BOS: begin
          BBRequest req = tagged IntSetHeader2BosReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_3_BOS: begin
          BBRequest req = tagged IntSetHeader3BosReqT {pkt: pkt};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_4_BOS: begin
          BBRequest req = tagged IntSetHeader4BosReqT {pkt: pkt};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_5_BOS: begin
          BBRequest req = tagged IntSetHeader5BosReqT {pkt: pkt};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_6_BOS: begin
          BBRequest req = tagged IntSetHeader6BosReqT {pkt: pkt};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_7_BOS: begin
          BBRequest req = tagged IntSetHeader7BosReqT {pkt: pkt};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntSetHeader0BosRspT {pkt: .pkt, int_switch_id_header$bos: .int_switch_id_header$bos}: begin
        meta.int_switch_id_header$bos = tagged Valid int_switch_id_header$bos;
        MetadataResponse rsp = tagged IntBosIntSetHeader0BosRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader1BosRspT {pkt: .pkt, int_ingress_port_id_header$bos: .int_ingress_port_id_header$bos}: begin
        meta.int_ingress_port_id_header$bos = tagged Valid int_ingress_port_id_header$bos;
        MetadataResponse rsp = tagged IntBosIntSetHeader1BosRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader2BosRspT {pkt: .pkt, int_hop_latency_header$bos: .int_hop_latency_header$bos}: begin
        meta.int_hop_latency_header$bos = tagged Valid int_hop_latency_header$bos;
        MetadataResponse rsp = tagged IntBosIntSetHeader2BosRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader3BosRspT {pkt: .pkt, int_q_occupancy_header$bos: .int_q_occupancy_header$bos}: begin
        meta.int_q_occupancy_header$bos = tagged Valid int_q_occupancy_header$bos;
        MetadataResponse rsp = tagged IntBosIntSetHeader3BosRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader4BosRspT {pkt: .pkt, int_ingress_tstamp_header$bos: .int_ingress_tstamp_header$bos}: begin
        meta.int_ingress_tstamp_header$bos = tagged Valid int_ingress_tstamp_header$bos;
        MetadataResponse rsp = tagged IntBosIntSetHeader4BosRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader5BosRspT {pkt: .pkt, int_egress_port_id_header$bos: .int_egress_port_id_header$bos}: begin
        meta.int_egress_port_id_header$bos = tagged Valid int_egress_port_id_header$bos;
        MetadataResponse rsp = tagged IntBosIntSetHeader5BosRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader6BosRspT {pkt: .pkt, int_q_congestion_header$bos: .int_q_congestion_header$bos}: begin
        meta.int_q_congestion_header$bos = tagged Valid int_q_congestion_header$bos;
        MetadataResponse rsp = tagged IntBosIntSetHeader6BosRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader7BosRspT {pkt: .pkt, int_egress_port_tx_utilization_header$bos: .int_egress_port_tx_utilization_header$bos}: begin
        meta.int_egress_port_tx_utilization_header$bos = tagged Valid int_egress_port_tx_utilization_header$bos;
        MetadataResponse rsp = tagged IntBosIntSetHeader7BosRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IntBosNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
endmodule

// ====== INT_INSERT ======

typedef struct {
  Bit#(6) padding;
  Bit#(1) int_metadata_i2e$source;
  Bit#(1) int_metadata_i2e$sink;
  Bit#(Bool) valid_int_header;
} IntInsertReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_INSERT,
  INT_TRANSIT,
  INT_SRC,
  INT_RESET
} IntInsertActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntInsertActionT _action;
  Bit#(32) runtime_switch_id;
  Bit#(8) runtime_hop_cnt;
  Bit#(5) runtime_ins_cnt;
  Bit#(4) runtime_ins_mask0003;
  Bit#(4) runtime_ins_mask0407;
  Bit#(16) runtime_ins_byte_cnt;
  Bit#(8) runtime_total_words;
} IntInsertRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(79)) matchtable_read_int_insert(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_int_insert(Bit#(9) msgtype, Bit#(79) data);
`endif
instance MatchTableSim#(111, 9, 79);
  function ActionValue#(Bit#(79)) matchtable_read(Bit#(111) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_int_insert(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(111) id, Bit#(9) key, Bit#(79) data);
    action
      matchtable_write_int_insert(key, data);
    endaction
  endfunction

endinstance
interface IntInsert;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIntInsert  (IntInsert);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(111, 256, SizeOf#(IntInsertReqT), SizeOf#(IntInsertRspT)) matchTable <- mkMatchTable("int_insert.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let int_metadata_i2e$source = fromMaybe(?, meta.int_metadata_i2e$source);
    let int_metadata_i2e$sink = fromMaybe(?, meta.int_metadata_i2e$sink);
    let i$n$t$_$h$e$a$d$e$r = fromMaybe(?, meta.i$n$t$_$h$e$a$d$e$r);
    IntInsertReqT req = IntInsertReqT {int_metadata_i2e$source: int_metadata_i2e$source,int_metadata_i2e$sink: int_metadata_i2e$sink,i$n$t$_$h$e$a$d$e$r: i$n$t$_$h$e$a$d$e$r};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntInsertRspT resp = unpack(data);
      case (resp._action) matches
        INT_TRANSIT: begin
          BBRequest req = tagged IntTransitReqT {pkt: pkt, int_header$ins_cnt: int_header$ins_cnt, runtime_switch_id: resp.runtime_switch_id};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INT_SRC: begin
          BBRequest req = tagged IntSrcReqT {pkt: pkt, runtime_total_words: resp.runtime_total_words, runtime_switch_id: resp.runtime_switch_id, runtime_ins_mask0003: resp.runtime_ins_mask0003, runtime_ins_byte_cnt: resp.runtime_ins_byte_cnt, runtime_ins_cnt: resp.runtime_ins_cnt, runtime_hop_cnt: resp.runtime_hop_cnt, runtime_ins_mask0407: resp.runtime_ins_mask0407};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        INT_RESET: begin
          BBRequest req = tagged IntResetReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntTransitRspT {pkt: .pkt, int_metadata$switch_id: .int_metadata$switch_id, int_metadata$gpe_int_hdr_len8: .int_metadata$gpe_int_hdr_len8}: begin
        meta.int_metadata$switch_id = tagged Valid int_metadata$switch_id;
        meta.int_metadata$gpe_int_hdr_len8 = tagged Valid int_metadata$gpe_int_hdr_len8;
        MetadataResponse rsp = tagged IntInsertIntTransitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSrcRspT {pkt: .pkt, int_metadata$gpe_int_hdr_len8: .int_metadata$gpe_int_hdr_len8, int_header$rsvd2: .int_header$rsvd2, int_header$ins_cnt: .int_header$ins_cnt, int_header$instruction_mask_0407: .int_header$instruction_mask_0407, int_header$total_hop_cnt: .int_header$total_hop_cnt, int_header$instruction_mask_1215: .int_header$instruction_mask_1215, int_header$rsvd1: .int_header$rsvd1, int_header$e: .int_header$e, int_header$instruction_mask_0811: .int_header$instruction_mask_0811, int_metadata$switch_id: .int_metadata$switch_id, int_header$rep: .int_header$rep, int_header$ver: .int_header$ver, int_header$max_hop_cnt: .int_header$max_hop_cnt, int_header$instruction_mask_0003: .int_header$instruction_mask_0003, int_metadata$insert_cnt: .int_metadata$insert_cnt, int_header$c: .int_header$c, int_metadata$insert_byte_cnt: .int_metadata$insert_byte_cnt}: begin
        meta.int_metadata$gpe_int_hdr_len8 = tagged Valid int_metadata$gpe_int_hdr_len8;
        meta.int_header$rsvd2 = tagged Valid int_header$rsvd2;
        meta.int_header$ins_cnt = tagged Valid int_header$ins_cnt;
        meta.int_header$instruction_mask_0407 = tagged Valid int_header$instruction_mask_0407;
        meta.int_header$total_hop_cnt = tagged Valid int_header$total_hop_cnt;
        meta.int_header$instruction_mask_1215 = tagged Valid int_header$instruction_mask_1215;
        meta.int_header$rsvd1 = tagged Valid int_header$rsvd1;
        meta.int_header$e = tagged Valid int_header$e;
        meta.int_header$instruction_mask_0811 = tagged Valid int_header$instruction_mask_0811;
        meta.int_metadata$switch_id = tagged Valid int_metadata$switch_id;
        meta.int_header$rep = tagged Valid int_header$rep;
        meta.int_header$ver = tagged Valid int_header$ver;
        meta.int_header$max_hop_cnt = tagged Valid int_header$max_hop_cnt;
        meta.int_header$instruction_mask_0003 = tagged Valid int_header$instruction_mask_0003;
        meta.int_metadata$insert_cnt = tagged Valid int_metadata$insert_cnt;
        meta.int_header$c = tagged Valid int_header$c;
        meta.int_metadata$insert_byte_cnt = tagged Valid int_metadata$insert_byte_cnt;
        MetadataResponse rsp = tagged IntInsertIntSrcRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntResetRspT {pkt: .pkt, int_metadata$switch_id: .int_metadata$switch_id, int_metadata$gpe_int_hdr_len8: .int_metadata$gpe_int_hdr_len8, int_metadata$insert_cnt: .int_metadata$insert_cnt, int_metadata$gpe_int_hdr_len: .int_metadata$gpe_int_hdr_len, int_metadata$insert_byte_cnt: .int_metadata$insert_byte_cnt, int_metadata$instruction_cnt: .int_metadata$instruction_cnt}: begin
        meta.int_metadata$switch_id = tagged Valid int_metadata$switch_id;
        meta.int_metadata$gpe_int_hdr_len8 = tagged Valid int_metadata$gpe_int_hdr_len8;
        meta.int_metadata$insert_cnt = tagged Valid int_metadata$insert_cnt;
        meta.int_metadata$gpe_int_hdr_len = tagged Valid int_metadata$gpe_int_hdr_len;
        meta.int_metadata$insert_byte_cnt = tagged Valid int_metadata$insert_byte_cnt;
        meta.int_metadata$instruction_cnt = tagged Valid int_metadata$instruction_cnt;
        MetadataResponse rsp = tagged IntInsertIntResetRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== INT_INST_0003 ======

typedef struct {
  Bit#(5) padding;
  Bit#(4) int_header$instruction_mask_0003;
} IntInst0003ReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_INST_0003,
  INT_SET_HEADER_0003_I0,
  INT_SET_HEADER_0003_I1,
  INT_SET_HEADER_0003_I2,
  INT_SET_HEADER_0003_I3,
  INT_SET_HEADER_0003_I4,
  INT_SET_HEADER_0003_I5,
  INT_SET_HEADER_0003_I6,
  INT_SET_HEADER_0003_I7,
  INT_SET_HEADER_0003_I8,
  INT_SET_HEADER_0003_I9,
  INT_SET_HEADER_0003_I10,
  INT_SET_HEADER_0003_I11,
  INT_SET_HEADER_0003_I12,
  INT_SET_HEADER_0003_I13,
  INT_SET_HEADER_0003_I14,
  INT_SET_HEADER_0003_I15
} IntInst0003ActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntInst0003ActionT _action;
} IntInst0003RspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(5)) matchtable_read_int_inst_0003(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_int_inst_0003(Bit#(9) msgtype, Bit#(5) data);
`endif
instance MatchTableSim#(105, 9, 5);
  function ActionValue#(Bit#(5)) matchtable_read(Bit#(105) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_int_inst_0003(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(105) id, Bit#(9) key, Bit#(5) data);
    action
      matchtable_write_int_inst_0003(key, data);
    endaction
  endfunction

endinstance
interface IntInst0003;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
  interface Client #(BBRequest, BBResponse) next_control_state_9;
  interface Client #(BBRequest, BBResponse) next_control_state_10;
  interface Client #(BBRequest, BBResponse) next_control_state_11;
  interface Client #(BBRequest, BBResponse) next_control_state_12;
  interface Client #(BBRequest, BBResponse) next_control_state_13;
  interface Client #(BBRequest, BBResponse) next_control_state_14;
  interface Client #(BBRequest, BBResponse) next_control_state_15;
endinterface
(* synthesize *)
module mkIntInst0003  (IntInst0003);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(16, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(16, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(105, 256, SizeOf#(IntInst0003ReqT), SizeOf#(IntInst0003RspT)) matchTable <- mkMatchTable("int_inst_0003.dat");
  Vector#(16, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(16) readyChannel = -1;
  for (Integer i=15; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let int_header$instruction_mask_0003 = fromMaybe(?, meta.int_header$instruction_mask_0003);
    IntInst0003ReqT req = IntInst0003ReqT {int_header$instruction_mask_0003: int_header$instruction_mask_0003};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntInst0003RspT resp = unpack(data);
      case (resp._action) matches
        INT_SET_HEADER_0003_I0: begin
          BBRequest req = tagged IntSetHeader0003I0ReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I1: begin
          BBRequest req = tagged IntSetHeader0003I1ReqT {pkt: pkt, intrinsic_metadata$enq_qdepth: intrinsic_metadata$enq_qdepth};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I2: begin
          BBRequest req = tagged IntSetHeader0003I2ReqT {pkt: pkt, intrinsic_metadata$deq_timedelta: intrinsic_metadata$deq_timedelta};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I3: begin
          BBRequest req = tagged IntSetHeader0003I3ReqT {pkt: pkt, intrinsic_metadata$deq_timedelta: intrinsic_metadata$deq_timedelta, intrinsic_metadata$enq_qdepth: intrinsic_metadata$enq_qdepth};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I4: begin
          BBRequest req = tagged IntSetHeader0003I4ReqT {pkt: pkt, ingress_metadata$ifindex: ingress_metadata$ifindex};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I5: begin
          BBRequest req = tagged IntSetHeader0003I5ReqT {pkt: pkt, intrinsic_metadata$enq_qdepth: intrinsic_metadata$enq_qdepth, ingress_metadata$ifindex: ingress_metadata$ifindex};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I6: begin
          BBRequest req = tagged IntSetHeader0003I6ReqT {pkt: pkt, intrinsic_metadata$deq_timedelta: intrinsic_metadata$deq_timedelta, ingress_metadata$ifindex: ingress_metadata$ifindex};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I7: begin
          BBRequest req = tagged IntSetHeader0003I7ReqT {pkt: pkt, intrinsic_metadata$deq_timedelta: intrinsic_metadata$deq_timedelta, intrinsic_metadata$enq_qdepth: intrinsic_metadata$enq_qdepth, ingress_metadata$ifindex: ingress_metadata$ifindex};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I8: begin
          BBRequest req = tagged IntSetHeader0003I8ReqT {pkt: pkt, int_metadata$switch_id: int_metadata$switch_id};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I9: begin
          BBRequest req = tagged IntSetHeader0003I9ReqT {pkt: pkt, int_metadata$switch_id: int_metadata$switch_id, intrinsic_metadata$enq_qdepth: intrinsic_metadata$enq_qdepth};
          bbReqFifo[9].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I10: begin
          BBRequest req = tagged IntSetHeader0003I10ReqT {pkt: pkt, intrinsic_metadata$deq_timedelta: intrinsic_metadata$deq_timedelta, int_metadata$switch_id: int_metadata$switch_id};
          bbReqFifo[10].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I11: begin
          BBRequest req = tagged IntSetHeader0003I11ReqT {pkt: pkt, intrinsic_metadata$deq_timedelta: intrinsic_metadata$deq_timedelta, intrinsic_metadata$enq_qdepth: intrinsic_metadata$enq_qdepth, int_metadata$switch_id: int_metadata$switch_id};
          bbReqFifo[11].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I12: begin
          BBRequest req = tagged IntSetHeader0003I12ReqT {pkt: pkt, int_metadata$switch_id: int_metadata$switch_id, ingress_metadata$ifindex: ingress_metadata$ifindex};
          bbReqFifo[12].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I13: begin
          BBRequest req = tagged IntSetHeader0003I13ReqT {pkt: pkt, int_metadata$switch_id: int_metadata$switch_id, intrinsic_metadata$enq_qdepth: intrinsic_metadata$enq_qdepth, ingress_metadata$ifindex: ingress_metadata$ifindex};
          bbReqFifo[13].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I14: begin
          BBRequest req = tagged IntSetHeader0003I14ReqT {pkt: pkt, intrinsic_metadata$deq_timedelta: intrinsic_metadata$deq_timedelta, ingress_metadata$ifindex: ingress_metadata$ifindex, int_metadata$switch_id: int_metadata$switch_id};
          bbReqFifo[14].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0003_I15: begin
          BBRequest req = tagged IntSetHeader0003I15ReqT {pkt: pkt, intrinsic_metadata$deq_timedelta: intrinsic_metadata$deq_timedelta, intrinsic_metadata$enq_qdepth: intrinsic_metadata$enq_qdepth, ingress_metadata$ifindex: ingress_metadata$ifindex, int_metadata$switch_id: int_metadata$switch_id};
          bbReqFifo[15].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntSetHeader0003I0RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I0RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I1RspT {pkt: .pkt, int_q_occupancy_header$q_occupancy0: .int_q_occupancy_header$q_occupancy0, int_q_occupancy_header$q_occupancy1: .int_q_occupancy_header$q_occupancy1}: begin
        meta.int_q_occupancy_header$q_occupancy0 = tagged Valid int_q_occupancy_header$q_occupancy0;
        meta.int_q_occupancy_header$q_occupancy1 = tagged Valid int_q_occupancy_header$q_occupancy1;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I2RspT {pkt: .pkt, int_hop_latency_header$hop_latency: .int_hop_latency_header$hop_latency}: begin
        meta.int_hop_latency_header$hop_latency = tagged Valid int_hop_latency_header$hop_latency;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I3RspT {pkt: .pkt, int_q_occupancy_header$q_occupancy0: .int_q_occupancy_header$q_occupancy0, int_hop_latency_header$hop_latency: .int_hop_latency_header$hop_latency, int_q_occupancy_header$q_occupancy1: .int_q_occupancy_header$q_occupancy1}: begin
        meta.int_q_occupancy_header$q_occupancy0 = tagged Valid int_q_occupancy_header$q_occupancy0;
        meta.int_hop_latency_header$hop_latency = tagged Valid int_hop_latency_header$hop_latency;
        meta.int_q_occupancy_header$q_occupancy1 = tagged Valid int_q_occupancy_header$q_occupancy1;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I4RspT {pkt: .pkt, int_ingress_port_id_header$ingress_port_id_1: .int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: .int_ingress_port_id_header$ingress_port_id_0}: begin
        meta.int_ingress_port_id_header$ingress_port_id_1 = tagged Valid int_ingress_port_id_header$ingress_port_id_1;
        meta.int_ingress_port_id_header$ingress_port_id_0 = tagged Valid int_ingress_port_id_header$ingress_port_id_0;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I5RspT {pkt: .pkt, int_ingress_port_id_header$ingress_port_id_1: .int_ingress_port_id_header$ingress_port_id_1, int_q_occupancy_header$q_occupancy0: .int_q_occupancy_header$q_occupancy0, int_ingress_port_id_header$ingress_port_id_0: .int_ingress_port_id_header$ingress_port_id_0, int_q_occupancy_header$q_occupancy1: .int_q_occupancy_header$q_occupancy1}: begin
        meta.int_ingress_port_id_header$ingress_port_id_1 = tagged Valid int_ingress_port_id_header$ingress_port_id_1;
        meta.int_q_occupancy_header$q_occupancy0 = tagged Valid int_q_occupancy_header$q_occupancy0;
        meta.int_ingress_port_id_header$ingress_port_id_0 = tagged Valid int_ingress_port_id_header$ingress_port_id_0;
        meta.int_q_occupancy_header$q_occupancy1 = tagged Valid int_q_occupancy_header$q_occupancy1;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I5RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I6RspT {pkt: .pkt, int_ingress_port_id_header$ingress_port_id_1: .int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: .int_ingress_port_id_header$ingress_port_id_0, int_hop_latency_header$hop_latency: .int_hop_latency_header$hop_latency}: begin
        meta.int_ingress_port_id_header$ingress_port_id_1 = tagged Valid int_ingress_port_id_header$ingress_port_id_1;
        meta.int_ingress_port_id_header$ingress_port_id_0 = tagged Valid int_ingress_port_id_header$ingress_port_id_0;
        meta.int_hop_latency_header$hop_latency = tagged Valid int_hop_latency_header$hop_latency;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I7RspT {pkt: .pkt, int_ingress_port_id_header$ingress_port_id_1: .int_ingress_port_id_header$ingress_port_id_1, int_q_occupancy_header$q_occupancy0: .int_q_occupancy_header$q_occupancy0, int_ingress_port_id_header$ingress_port_id_0: .int_ingress_port_id_header$ingress_port_id_0, int_hop_latency_header$hop_latency: .int_hop_latency_header$hop_latency, int_q_occupancy_header$q_occupancy1: .int_q_occupancy_header$q_occupancy1}: begin
        meta.int_ingress_port_id_header$ingress_port_id_1 = tagged Valid int_ingress_port_id_header$ingress_port_id_1;
        meta.int_q_occupancy_header$q_occupancy0 = tagged Valid int_q_occupancy_header$q_occupancy0;
        meta.int_ingress_port_id_header$ingress_port_id_0 = tagged Valid int_ingress_port_id_header$ingress_port_id_0;
        meta.int_hop_latency_header$hop_latency = tagged Valid int_hop_latency_header$hop_latency;
        meta.int_q_occupancy_header$q_occupancy1 = tagged Valid int_q_occupancy_header$q_occupancy1;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I7RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I8RspT {pkt: .pkt, int_switch_id_header$switch_id: .int_switch_id_header$switch_id}: begin
        meta.int_switch_id_header$switch_id = tagged Valid int_switch_id_header$switch_id;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I8RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I9RspT {pkt: .pkt, int_q_occupancy_header$q_occupancy0: .int_q_occupancy_header$q_occupancy0, int_switch_id_header$switch_id: .int_switch_id_header$switch_id, int_q_occupancy_header$q_occupancy1: .int_q_occupancy_header$q_occupancy1}: begin
        meta.int_q_occupancy_header$q_occupancy0 = tagged Valid int_q_occupancy_header$q_occupancy0;
        meta.int_switch_id_header$switch_id = tagged Valid int_switch_id_header$switch_id;
        meta.int_q_occupancy_header$q_occupancy1 = tagged Valid int_q_occupancy_header$q_occupancy1;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I9RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I10RspT {pkt: .pkt, int_switch_id_header$switch_id: .int_switch_id_header$switch_id, int_hop_latency_header$hop_latency: .int_hop_latency_header$hop_latency}: begin
        meta.int_switch_id_header$switch_id = tagged Valid int_switch_id_header$switch_id;
        meta.int_hop_latency_header$hop_latency = tagged Valid int_hop_latency_header$hop_latency;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I10RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I11RspT {pkt: .pkt, int_switch_id_header$switch_id: .int_switch_id_header$switch_id, int_q_occupancy_header$q_occupancy0: .int_q_occupancy_header$q_occupancy0, int_hop_latency_header$hop_latency: .int_hop_latency_header$hop_latency, int_q_occupancy_header$q_occupancy1: .int_q_occupancy_header$q_occupancy1}: begin
        meta.int_switch_id_header$switch_id = tagged Valid int_switch_id_header$switch_id;
        meta.int_q_occupancy_header$q_occupancy0 = tagged Valid int_q_occupancy_header$q_occupancy0;
        meta.int_hop_latency_header$hop_latency = tagged Valid int_hop_latency_header$hop_latency;
        meta.int_q_occupancy_header$q_occupancy1 = tagged Valid int_q_occupancy_header$q_occupancy1;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I11RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I12RspT {pkt: .pkt, int_ingress_port_id_header$ingress_port_id_1: .int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: .int_ingress_port_id_header$ingress_port_id_0, int_switch_id_header$switch_id: .int_switch_id_header$switch_id}: begin
        meta.int_ingress_port_id_header$ingress_port_id_1 = tagged Valid int_ingress_port_id_header$ingress_port_id_1;
        meta.int_ingress_port_id_header$ingress_port_id_0 = tagged Valid int_ingress_port_id_header$ingress_port_id_0;
        meta.int_switch_id_header$switch_id = tagged Valid int_switch_id_header$switch_id;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I12RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I13RspT {pkt: .pkt, int_ingress_port_id_header$ingress_port_id_1: .int_ingress_port_id_header$ingress_port_id_1, int_q_occupancy_header$q_occupancy0: .int_q_occupancy_header$q_occupancy0, int_ingress_port_id_header$ingress_port_id_0: .int_ingress_port_id_header$ingress_port_id_0, int_switch_id_header$switch_id: .int_switch_id_header$switch_id, int_q_occupancy_header$q_occupancy1: .int_q_occupancy_header$q_occupancy1}: begin
        meta.int_ingress_port_id_header$ingress_port_id_1 = tagged Valid int_ingress_port_id_header$ingress_port_id_1;
        meta.int_q_occupancy_header$q_occupancy0 = tagged Valid int_q_occupancy_header$q_occupancy0;
        meta.int_ingress_port_id_header$ingress_port_id_0 = tagged Valid int_ingress_port_id_header$ingress_port_id_0;
        meta.int_switch_id_header$switch_id = tagged Valid int_switch_id_header$switch_id;
        meta.int_q_occupancy_header$q_occupancy1 = tagged Valid int_q_occupancy_header$q_occupancy1;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I13RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I14RspT {pkt: .pkt, int_ingress_port_id_header$ingress_port_id_1: .int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: .int_ingress_port_id_header$ingress_port_id_0, int_switch_id_header$switch_id: .int_switch_id_header$switch_id, int_hop_latency_header$hop_latency: .int_hop_latency_header$hop_latency}: begin
        meta.int_ingress_port_id_header$ingress_port_id_1 = tagged Valid int_ingress_port_id_header$ingress_port_id_1;
        meta.int_ingress_port_id_header$ingress_port_id_0 = tagged Valid int_ingress_port_id_header$ingress_port_id_0;
        meta.int_switch_id_header$switch_id = tagged Valid int_switch_id_header$switch_id;
        meta.int_hop_latency_header$hop_latency = tagged Valid int_hop_latency_header$hop_latency;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I14RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0003I15RspT {pkt: .pkt, int_q_occupancy_header$q_occupancy0: .int_q_occupancy_header$q_occupancy0, int_switch_id_header$switch_id: .int_switch_id_header$switch_id, int_hop_latency_header$hop_latency: .int_hop_latency_header$hop_latency, int_ingress_port_id_header$ingress_port_id_1: .int_ingress_port_id_header$ingress_port_id_1, int_ingress_port_id_header$ingress_port_id_0: .int_ingress_port_id_header$ingress_port_id_0, int_q_occupancy_header$q_occupancy1: .int_q_occupancy_header$q_occupancy1}: begin
        meta.int_q_occupancy_header$q_occupancy0 = tagged Valid int_q_occupancy_header$q_occupancy0;
        meta.int_switch_id_header$switch_id = tagged Valid int_switch_id_header$switch_id;
        meta.int_hop_latency_header$hop_latency = tagged Valid int_hop_latency_header$hop_latency;
        meta.int_ingress_port_id_header$ingress_port_id_1 = tagged Valid int_ingress_port_id_header$ingress_port_id_1;
        meta.int_ingress_port_id_header$ingress_port_id_0 = tagged Valid int_ingress_port_id_header$ingress_port_id_0;
        meta.int_q_occupancy_header$q_occupancy1 = tagged Valid int_q_occupancy_header$q_occupancy1;
        MetadataResponse rsp = tagged IntInst0003IntSetHeader0003I15RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
  interface next_control_state_9 = toClient(bbReqFifo[9], bbRspFifo[9]);
  interface next_control_state_10 = toClient(bbReqFifo[10], bbRspFifo[10]);
  interface next_control_state_11 = toClient(bbReqFifo[11], bbRspFifo[11]);
  interface next_control_state_12 = toClient(bbReqFifo[12], bbRspFifo[12]);
  interface next_control_state_13 = toClient(bbReqFifo[13], bbRspFifo[13]);
  interface next_control_state_14 = toClient(bbReqFifo[14], bbRspFifo[14]);
  interface next_control_state_15 = toClient(bbReqFifo[15], bbRspFifo[15]);
endmodule

// ====== INT_INST_0407 ======

typedef struct {
  Bit#(5) padding;
  Bit#(4) int_header$instruction_mask_0407;
} IntInst0407ReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_INST_0407,
  INT_SET_HEADER_0407_I0,
  INT_SET_HEADER_0407_I1,
  INT_SET_HEADER_0407_I2,
  INT_SET_HEADER_0407_I3,
  INT_SET_HEADER_0407_I4,
  INT_SET_HEADER_0407_I5,
  INT_SET_HEADER_0407_I6,
  INT_SET_HEADER_0407_I7,
  INT_SET_HEADER_0407_I8,
  INT_SET_HEADER_0407_I9,
  INT_SET_HEADER_0407_I10,
  INT_SET_HEADER_0407_I11,
  INT_SET_HEADER_0407_I12,
  INT_SET_HEADER_0407_I13,
  INT_SET_HEADER_0407_I14,
  INT_SET_HEADER_0407_I15,
  NOP
} IntInst0407ActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntInst0407ActionT _action;
} IntInst0407RspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(5)) matchtable_read_int_inst_0407(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_int_inst_0407(Bit#(9) msgtype, Bit#(5) data);
`endif
instance MatchTableSim#(106, 9, 5);
  function ActionValue#(Bit#(5)) matchtable_read(Bit#(106) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_int_inst_0407(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(106) id, Bit#(9) key, Bit#(5) data);
    action
      matchtable_write_int_inst_0407(key, data);
    endaction
  endfunction

endinstance
interface IntInst0407;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
  interface Client #(BBRequest, BBResponse) next_control_state_9;
  interface Client #(BBRequest, BBResponse) next_control_state_10;
  interface Client #(BBRequest, BBResponse) next_control_state_11;
  interface Client #(BBRequest, BBResponse) next_control_state_12;
  interface Client #(BBRequest, BBResponse) next_control_state_13;
  interface Client #(BBRequest, BBResponse) next_control_state_14;
  interface Client #(BBRequest, BBResponse) next_control_state_15;
  interface Client #(BBRequest, BBResponse) next_control_state_16;
endinterface
(* synthesize *)
module mkIntInst0407  (IntInst0407);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(17, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(17, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(106, 256, SizeOf#(IntInst0407ReqT), SizeOf#(IntInst0407RspT)) matchTable <- mkMatchTable("int_inst_0407.dat");
  Vector#(17, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(17) readyChannel = -1;
  for (Integer i=16; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let int_header$instruction_mask_0407 = fromMaybe(?, meta.int_header$instruction_mask_0407);
    IntInst0407ReqT req = IntInst0407ReqT {int_header$instruction_mask_0407: int_header$instruction_mask_0407};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntInst0407RspT resp = unpack(data);
      case (resp._action) matches
        INT_SET_HEADER_0407_I0: begin
          BBRequest req = tagged IntSetHeader0407I0ReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I1: begin
          BBRequest req = tagged IntSetHeader0407I1ReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I2: begin
          BBRequest req = tagged IntSetHeader0407I2ReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I3: begin
          BBRequest req = tagged IntSetHeader0407I3ReqT {pkt: pkt};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I4: begin
          BBRequest req = tagged IntSetHeader0407I4ReqT {pkt: pkt, standard_metadata$egress_port: standard_metadata$egress_port};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I5: begin
          BBRequest req = tagged IntSetHeader0407I5ReqT {pkt: pkt, standard_metadata$egress_port: standard_metadata$egress_port};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I6: begin
          BBRequest req = tagged IntSetHeader0407I6ReqT {pkt: pkt, standard_metadata$egress_port: standard_metadata$egress_port};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I7: begin
          BBRequest req = tagged IntSetHeader0407I7ReqT {pkt: pkt, standard_metadata$egress_port: standard_metadata$egress_port};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I8: begin
          BBRequest req = tagged IntSetHeader0407I8ReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I9: begin
          BBRequest req = tagged IntSetHeader0407I9ReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp};
          bbReqFifo[9].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I10: begin
          BBRequest req = tagged IntSetHeader0407I10ReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp};
          bbReqFifo[10].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I11: begin
          BBRequest req = tagged IntSetHeader0407I11ReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp};
          bbReqFifo[11].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I12: begin
          BBRequest req = tagged IntSetHeader0407I12ReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp, standard_metadata$egress_port: standard_metadata$egress_port};
          bbReqFifo[12].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I13: begin
          BBRequest req = tagged IntSetHeader0407I13ReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp, standard_metadata$egress_port: standard_metadata$egress_port};
          bbReqFifo[13].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I14: begin
          BBRequest req = tagged IntSetHeader0407I14ReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp, standard_metadata$egress_port: standard_metadata$egress_port};
          bbReqFifo[14].enq(req); //FIXME: replace with RXTX.
        end
        INT_SET_HEADER_0407_I15: begin
          BBRequest req = tagged IntSetHeader0407I15ReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp, standard_metadata$egress_port: standard_metadata$egress_port};
          bbReqFifo[15].enq(req); //FIXME: replace with RXTX.
        end
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[16].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntSetHeader0407I0RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I0RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I1RspT {pkt: .pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: .int_egress_port_tx_utilization_header$egress_port_tx_utilization}: begin
        meta.int_egress_port_tx_utilization_header$egress_port_tx_utilization = tagged Valid int_egress_port_tx_utilization_header$egress_port_tx_utilization;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I2RspT {pkt: .pkt, int_q_congestion_header$q_congestion: .int_q_congestion_header$q_congestion}: begin
        meta.int_q_congestion_header$q_congestion = tagged Valid int_q_congestion_header$q_congestion;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I3RspT {pkt: .pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: .int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_q_congestion_header$q_congestion: .int_q_congestion_header$q_congestion}: begin
        meta.int_egress_port_tx_utilization_header$egress_port_tx_utilization = tagged Valid int_egress_port_tx_utilization_header$egress_port_tx_utilization;
        meta.int_q_congestion_header$q_congestion = tagged Valid int_q_congestion_header$q_congestion;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I4RspT {pkt: .pkt, int_egress_port_id_header$egress_port_id: .int_egress_port_id_header$egress_port_id}: begin
        meta.int_egress_port_id_header$egress_port_id = tagged Valid int_egress_port_id_header$egress_port_id;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I5RspT {pkt: .pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: .int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_egress_port_id_header$egress_port_id: .int_egress_port_id_header$egress_port_id}: begin
        meta.int_egress_port_tx_utilization_header$egress_port_tx_utilization = tagged Valid int_egress_port_tx_utilization_header$egress_port_tx_utilization;
        meta.int_egress_port_id_header$egress_port_id = tagged Valid int_egress_port_id_header$egress_port_id;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I5RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I6RspT {pkt: .pkt, int_q_congestion_header$q_congestion: .int_q_congestion_header$q_congestion, int_egress_port_id_header$egress_port_id: .int_egress_port_id_header$egress_port_id}: begin
        meta.int_q_congestion_header$q_congestion = tagged Valid int_q_congestion_header$q_congestion;
        meta.int_egress_port_id_header$egress_port_id = tagged Valid int_egress_port_id_header$egress_port_id;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I7RspT {pkt: .pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: .int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_egress_port_id_header$egress_port_id: .int_egress_port_id_header$egress_port_id, int_q_congestion_header$q_congestion: .int_q_congestion_header$q_congestion}: begin
        meta.int_egress_port_tx_utilization_header$egress_port_tx_utilization = tagged Valid int_egress_port_tx_utilization_header$egress_port_tx_utilization;
        meta.int_egress_port_id_header$egress_port_id = tagged Valid int_egress_port_id_header$egress_port_id;
        meta.int_q_congestion_header$q_congestion = tagged Valid int_q_congestion_header$q_congestion;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I7RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I8RspT {pkt: .pkt, int_ingress_tstamp_header$ingress_tstamp: .int_ingress_tstamp_header$ingress_tstamp}: begin
        meta.int_ingress_tstamp_header$ingress_tstamp = tagged Valid int_ingress_tstamp_header$ingress_tstamp;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I8RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I9RspT {pkt: .pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: .int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_ingress_tstamp_header$ingress_tstamp: .int_ingress_tstamp_header$ingress_tstamp}: begin
        meta.int_egress_port_tx_utilization_header$egress_port_tx_utilization = tagged Valid int_egress_port_tx_utilization_header$egress_port_tx_utilization;
        meta.int_ingress_tstamp_header$ingress_tstamp = tagged Valid int_ingress_tstamp_header$ingress_tstamp;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I9RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I10RspT {pkt: .pkt, int_q_congestion_header$q_congestion: .int_q_congestion_header$q_congestion, int_ingress_tstamp_header$ingress_tstamp: .int_ingress_tstamp_header$ingress_tstamp}: begin
        meta.int_q_congestion_header$q_congestion = tagged Valid int_q_congestion_header$q_congestion;
        meta.int_ingress_tstamp_header$ingress_tstamp = tagged Valid int_ingress_tstamp_header$ingress_tstamp;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I10RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I11RspT {pkt: .pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: .int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_q_congestion_header$q_congestion: .int_q_congestion_header$q_congestion, int_ingress_tstamp_header$ingress_tstamp: .int_ingress_tstamp_header$ingress_tstamp}: begin
        meta.int_egress_port_tx_utilization_header$egress_port_tx_utilization = tagged Valid int_egress_port_tx_utilization_header$egress_port_tx_utilization;
        meta.int_q_congestion_header$q_congestion = tagged Valid int_q_congestion_header$q_congestion;
        meta.int_ingress_tstamp_header$ingress_tstamp = tagged Valid int_ingress_tstamp_header$ingress_tstamp;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I11RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I12RspT {pkt: .pkt, int_egress_port_id_header$egress_port_id: .int_egress_port_id_header$egress_port_id, int_ingress_tstamp_header$ingress_tstamp: .int_ingress_tstamp_header$ingress_tstamp}: begin
        meta.int_egress_port_id_header$egress_port_id = tagged Valid int_egress_port_id_header$egress_port_id;
        meta.int_ingress_tstamp_header$ingress_tstamp = tagged Valid int_ingress_tstamp_header$ingress_tstamp;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I12RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I13RspT {pkt: .pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: .int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_egress_port_id_header$egress_port_id: .int_egress_port_id_header$egress_port_id, int_ingress_tstamp_header$ingress_tstamp: .int_ingress_tstamp_header$ingress_tstamp}: begin
        meta.int_egress_port_tx_utilization_header$egress_port_tx_utilization = tagged Valid int_egress_port_tx_utilization_header$egress_port_tx_utilization;
        meta.int_egress_port_id_header$egress_port_id = tagged Valid int_egress_port_id_header$egress_port_id;
        meta.int_ingress_tstamp_header$ingress_tstamp = tagged Valid int_ingress_tstamp_header$ingress_tstamp;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I13RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I14RspT {pkt: .pkt, int_q_congestion_header$q_congestion: .int_q_congestion_header$q_congestion, int_egress_port_id_header$egress_port_id: .int_egress_port_id_header$egress_port_id, int_ingress_tstamp_header$ingress_tstamp: .int_ingress_tstamp_header$ingress_tstamp}: begin
        meta.int_q_congestion_header$q_congestion = tagged Valid int_q_congestion_header$q_congestion;
        meta.int_egress_port_id_header$egress_port_id = tagged Valid int_egress_port_id_header$egress_port_id;
        meta.int_ingress_tstamp_header$ingress_tstamp = tagged Valid int_ingress_tstamp_header$ingress_tstamp;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I14RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntSetHeader0407I15RspT {pkt: .pkt, int_egress_port_tx_utilization_header$egress_port_tx_utilization: .int_egress_port_tx_utilization_header$egress_port_tx_utilization, int_egress_port_id_header$egress_port_id: .int_egress_port_id_header$egress_port_id, int_q_congestion_header$q_congestion: .int_q_congestion_header$q_congestion, int_ingress_tstamp_header$ingress_tstamp: .int_ingress_tstamp_header$ingress_tstamp}: begin
        meta.int_egress_port_tx_utilization_header$egress_port_tx_utilization = tagged Valid int_egress_port_tx_utilization_header$egress_port_tx_utilization;
        meta.int_egress_port_id_header$egress_port_id = tagged Valid int_egress_port_id_header$egress_port_id;
        meta.int_q_congestion_header$q_congestion = tagged Valid int_q_congestion_header$q_congestion;
        meta.int_ingress_tstamp_header$ingress_tstamp = tagged Valid int_ingress_tstamp_header$ingress_tstamp;
        MetadataResponse rsp = tagged IntInst0407IntSetHeader0407I15RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IntInst0407NopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
  interface next_control_state_9 = toClient(bbReqFifo[9], bbRspFifo[9]);
  interface next_control_state_10 = toClient(bbReqFifo[10], bbRspFifo[10]);
  interface next_control_state_11 = toClient(bbReqFifo[11], bbRspFifo[11]);
  interface next_control_state_12 = toClient(bbReqFifo[12], bbRspFifo[12]);
  interface next_control_state_13 = toClient(bbReqFifo[13], bbRspFifo[13]);
  interface next_control_state_14 = toClient(bbReqFifo[14], bbRspFifo[14]);
  interface next_control_state_15 = toClient(bbReqFifo[15], bbRspFifo[15]);
  interface next_control_state_16 = toClient(bbReqFifo[16], bbRspFifo[16]);
endmodule

// ====== INT_INST_0811 ======

typedef struct {
  Bit#(5) padding;
  Bit#(4) int_header$instruction_mask_0811;
} IntInst0811ReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_INST_0811,
  NOP
} IntInst0811ActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntInst0811ActionT _action;
} IntInst0811RspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_int_inst_0811(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_int_inst_0811(Bit#(9) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(107, 9, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(107) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_int_inst_0811(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(107) id, Bit#(9) key, Bit#(1) data);
    action
      matchtable_write_int_inst_0811(key, data);
    endaction
  endfunction

endinstance
interface IntInst0811;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkIntInst0811  (IntInst0811);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(107, 256, SizeOf#(IntInst0811ReqT), SizeOf#(IntInst0811RspT)) matchTable <- mkMatchTable("int_inst_0811.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let int_header$instruction_mask_0811 = fromMaybe(?, meta.int_header$instruction_mask_0811);
    IntInst0811ReqT req = IntInst0811ReqT {int_header$instruction_mask_0811: int_header$instruction_mask_0811};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntInst0811RspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IntInst0811NopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== INT_INST_1215 ======

typedef struct {
  Bit#(5) padding;
  Bit#(4) int_header$instruction_mask_1215;
} IntInst1215ReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_INST_1215,
  NOP
} IntInst1215ActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntInst1215ActionT _action;
} IntInst1215RspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(1)) matchtable_read_int_inst_1215(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_int_inst_1215(Bit#(9) msgtype, Bit#(1) data);
`endif
instance MatchTableSim#(108, 9, 1);
  function ActionValue#(Bit#(1)) matchtable_read(Bit#(108) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_int_inst_1215(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(108) id, Bit#(9) key, Bit#(1) data);
    action
      matchtable_write_int_inst_1215(key, data);
    endaction
  endfunction

endinstance
interface IntInst1215;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkIntInst1215  (IntInst1215);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(108, 256, SizeOf#(IntInst1215ReqT), SizeOf#(IntInst1215RspT)) matchTable <- mkMatchTable("int_inst_1215.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let int_header$instruction_mask_1215 = fromMaybe(?, meta.int_header$instruction_mask_1215);
    IntInst1215ReqT req = IntInst1215ReqT {int_header$instruction_mask_1215: int_header$instruction_mask_1215};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntInst1215RspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IntInst1215NopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== INT_META_HEADER_UPDATE ======

typedef struct {
  Bit#(1) padding;
  Bit#(8) int_metadata$insert_cnt;
} IntMetaHeaderUpdateReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_META_HEADER_UPDATE,
  INT_SET_E_BIT,
  INT_UPDATE_TOTAL_HOP_CNT
} IntMetaHeaderUpdateActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntMetaHeaderUpdateActionT _action;
} IntMetaHeaderUpdateRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_int_meta_header_update(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_int_meta_header_update(Bit#(9) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(110, 9, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(110) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_int_meta_header_update(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(110) id, Bit#(9) key, Bit#(2) data);
    action
      matchtable_write_int_meta_header_update(key, data);
    endaction
  endfunction

endinstance
interface IntMetaHeaderUpdate;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkIntMetaHeaderUpdate  (IntMetaHeaderUpdate);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(110, 256, SizeOf#(IntMetaHeaderUpdateReqT), SizeOf#(IntMetaHeaderUpdateRspT)) matchTable <- mkMatchTable("int_meta_header_update.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let int_metadata$insert_cnt = fromMaybe(?, meta.int_metadata$insert_cnt);
    IntMetaHeaderUpdateReqT req = IntMetaHeaderUpdateReqT {int_metadata$insert_cnt: int_metadata$insert_cnt};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntMetaHeaderUpdateRspT resp = unpack(data);
      case (resp._action) matches
        INT_SET_E_BIT: begin
          BBRequest req = tagged IntSetEBitReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INT_UPDATE_TOTAL_HOP_CNT: begin
          BBRequest req = tagged IntUpdateTotalHopCntReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntSetEBitRspT {pkt: .pkt, int_header$e: .int_header$e}: begin
        meta.int_header$e = tagged Valid int_header$e;
        MetadataResponse rsp = tagged IntMetaHeaderUpdateIntSetEBitRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntUpdateTotalHopCntRspT {pkt: .pkt, int_header$total_hop_cnt: .int_header$total_hop_cnt}: begin
        meta.int_header$total_hop_cnt = tagged Valid int_header$total_hop_cnt;
        MetadataResponse rsp = tagged IntMetaHeaderUpdateIntUpdateTotalHopCntRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== INT_OUTER_ENCAP ======

typedef struct {
  Bit#(1) padding;
  Bit#(Bool) valid_ipv4;
  Bit#(Bool) valid_vxlan_gpe;
  Bit#(1) int_metadata_i2e$source;
  Bit#(5) tunnel_metadata$egress_tunnel_type;
} IntOuterEncapReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_INT_OUTER_ENCAP,
  INT_UPDATE_VXLAN_GPE_IPV4,
  INT_ADD_UPDATE_VXLAN_GPE_IPV4,
  NOP
} IntOuterEncapActionT deriving (Bits, Eq, FShow);
typedef struct {
  IntOuterEncapActionT _action;
} IntOuterEncapRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_int_outer_encap(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_int_outer_encap(Bit#(9) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(112, 9, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(112) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_int_outer_encap(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(112) id, Bit#(9) key, Bit#(2) data);
    action
      matchtable_write_int_outer_encap(key, data);
    endaction
  endfunction

endinstance
interface IntOuterEncap;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkIntOuterEncap  (IntOuterEncap);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(112, 256, SizeOf#(IntOuterEncapReqT), SizeOf#(IntOuterEncapRspT)) matchTable <- mkMatchTable("int_outer_encap.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let v$x$l$a$n$_$g$p$e = fromMaybe(?, meta.v$x$l$a$n$_$g$p$e);
    let int_metadata_i2e$source = fromMaybe(?, meta.int_metadata_i2e$source);
    let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
    IntOuterEncapReqT req = IntOuterEncapReqT {i$p$v$4: i$p$v$4,v$x$l$a$n$_$g$p$e: v$x$l$a$n$_$g$p$e,int_metadata_i2e$source: int_metadata_i2e$source,tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      IntOuterEncapRspT resp = unpack(data);
      case (resp._action) matches
        INT_UPDATE_VXLAN_GPE_IPV4: begin
          BBRequest req = tagged IntUpdateVxlanGpeIpv4ReqT {pkt: pkt, int_metadata$gpe_int_hdr_len8: int_metadata$gpe_int_hdr_len8, int_metadata$insert_byte_cnt: int_metadata$insert_byte_cnt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INT_ADD_UPDATE_VXLAN_GPE_IPV4: begin
          BBRequest req = tagged IntAddUpdateVxlanGpeIpv4ReqT {pkt: pkt, int_metadata$gpe_int_hdr_len8: int_metadata$gpe_int_hdr_len8, int_metadata$insert_byte_cnt: int_metadata$insert_byte_cnt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged IntUpdateVxlanGpeIpv4RspT {pkt: .pkt, vxlan_gpe_int_header$len: .vxlan_gpe_int_header$len, udp$length_: .udp$length_, ipv4$totalLen: .ipv4$totalLen}: begin
        meta.vxlan_gpe_int_header$len = tagged Valid vxlan_gpe_int_header$len;
        meta.udp$length_ = tagged Valid udp$length_;
        meta.ipv4$totalLen = tagged Valid ipv4$totalLen;
        MetadataResponse rsp = tagged IntOuterEncapIntUpdateVxlanGpeIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged IntAddUpdateVxlanGpeIpv4RspT {pkt: .pkt, vxlan_gpe$next_proto: .vxlan_gpe$next_proto, vxlan_gpe_int_header$len: .vxlan_gpe_int_header$len, vxlan_gpe_int_header$next_proto: .vxlan_gpe_int_header$next_proto, vxlan_gpe_int_header$int_type: .vxlan_gpe_int_header$int_type, udp$length_: .udp$length_, ipv4$totalLen: .ipv4$totalLen}: begin
        meta.vxlan_gpe$next_proto = tagged Valid vxlan_gpe$next_proto;
        meta.vxlan_gpe_int_header$len = tagged Valid vxlan_gpe_int_header$len;
        meta.vxlan_gpe_int_header$next_proto = tagged Valid vxlan_gpe_int_header$next_proto;
        meta.vxlan_gpe_int_header$int_type = tagged Valid vxlan_gpe_int_header$int_type;
        meta.udp$length_ = tagged Valid udp$length_;
        meta.ipv4$totalLen = tagged Valid ipv4$totalLen;
        MetadataResponse rsp = tagged IntOuterEncapIntAddUpdateVxlanGpeIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged IntOuterEncapNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== L3_REWRITE ======

typedef struct {
  Bit#(8) padding;
  Bit#(Bool) valid_ipv4;
  Bit#(Bool) valid_ipv6;
  Bit#(Bool) valid_mpls0;
  Bit#(32) ipv4$dstAddr;
  Bit#(128) ipv6$dstAddr;
} L3RewriteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_L3_REWRITE,
  NOP,
  IPV4_UNICAST_REWRITE,
  IPV4_MULTICAST_REWRITE,
  IPV6_UNICAST_REWRITE,
  IPV6_MULTICAST_REWRITE,
  MPLS_REWRITE
} L3RewriteActionT deriving (Bits, Eq, FShow);
typedef struct {
  L3RewriteActionT _action;
} L3RewriteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(3)) matchtable_read_l3_rewrite(Bit#(171) msgtype);
import "BDPI" function Action matchtable_write_l3_rewrite(Bit#(171) msgtype, Bit#(3) data);
`endif
instance MatchTableSim#(84, 171, 3);
  function ActionValue#(Bit#(3)) matchtable_read(Bit#(84) id, Bit#(171) key);
    actionvalue
      let v <- matchtable_read_l3_rewrite(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(84) id, Bit#(171) key, Bit#(3) data);
    action
      matchtable_write_l3_rewrite(key, data);
    endaction
  endfunction

endinstance
interface L3Rewrite;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
endinterface
(* synthesize *)
module mkL3Rewrite  (L3Rewrite);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(6, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(6, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(84, 256, SizeOf#(L3RewriteReqT), SizeOf#(L3RewriteRspT)) matchTable <- mkMatchTable("l3_rewrite.dat");
  Vector#(6, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(6) readyChannel = -1;
  for (Integer i=5; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let i$p$v$6 = fromMaybe(?, meta.i$p$v$6);
    let m$p$l$s$$0$ = fromMaybe(?, meta.m$p$l$s$$0$);
    let ipv4$dstAddr = fromMaybe(?, meta.ipv4$dstAddr);
    let ipv6$dstAddr = fromMaybe(?, meta.ipv6$dstAddr);
    L3RewriteReqT req = L3RewriteReqT {i$p$v$4: i$p$v$4,i$p$v$6: i$p$v$6,m$p$l$s$$0$: m$p$l$s$$0$,ipv4$dstAddr: ipv4$dstAddr,ipv6$dstAddr: ipv6$dstAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      L3RewriteRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_UNICAST_REWRITE: begin
          BBRequest req = tagged Ipv4UnicastRewriteReqT {pkt: pkt, egress_metadata$mac_da: egress_metadata$mac_da};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_MULTICAST_REWRITE: begin
          BBRequest req = tagged Ipv4MulticastRewriteReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_UNICAST_REWRITE: begin
          BBRequest req = tagged Ipv6UnicastRewriteReqT {pkt: pkt, egress_metadata$mac_da: egress_metadata$mac_da};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_MULTICAST_REWRITE: begin
          BBRequest req = tagged Ipv6MulticastRewriteReqT {pkt: pkt};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        MPLS_REWRITE: begin
          BBRequest req = tagged MplsRewriteReqT {pkt: pkt, egress_metadata$mac_da: egress_metadata$mac_da};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged L3RewriteNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4UnicastRewriteRspT {pkt: .pkt, ipv4$ttl: .ipv4$ttl, ethernet$dstAddr: .ethernet$dstAddr}: begin
        meta.ipv4$ttl = tagged Valid ipv4$ttl;
        meta.ethernet$dstAddr = tagged Valid ethernet$dstAddr;
        MetadataResponse rsp = tagged L3RewriteIpv4UnicastRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4MulticastRewriteRspT {pkt: .pkt, ipv4$ttl: .ipv4$ttl}: begin
        meta.ipv4$ttl = tagged Valid ipv4$ttl;
        MetadataResponse rsp = tagged L3RewriteIpv4MulticastRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6UnicastRewriteRspT {pkt: .pkt, ipv6$hopLimit: .ipv6$hopLimit, ethernet$dstAddr: .ethernet$dstAddr}: begin
        meta.ipv6$hopLimit = tagged Valid ipv6$hopLimit;
        meta.ethernet$dstAddr = tagged Valid ethernet$dstAddr;
        MetadataResponse rsp = tagged L3RewriteIpv6UnicastRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6MulticastRewriteRspT {pkt: .pkt, ipv6$hopLimit: .ipv6$hopLimit}: begin
        meta.ipv6$hopLimit = tagged Valid ipv6$hopLimit;
        MetadataResponse rsp = tagged L3RewriteIpv6MulticastRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MplsRewriteRspT {pkt: .pkt, ethernet$dstAddr: .ethernet$dstAddr, mpls0$ttl: .mpls0$ttl}: begin
        meta.ethernet$dstAddr = tagged Valid ethernet$dstAddr;
        meta.mpls0$ttl = tagged Valid mpls0$ttl;
        MetadataResponse rsp = tagged L3RewriteMplsRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
endmodule

// ====== MIRROR ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) i2e_metadata$mirror_session_id;
} MirrorReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_MIRROR,
  NOP,
  SET_MIRROR_NHOP,
  SET_MIRROR_BD,
  SFLOW_PKT_TO_CPU
} MirrorActionT deriving (Bits, Eq, FShow);
typedef struct {
  MirrorActionT _action;
  Bit#(16) runtime_nhop_idx;
  Bit#(16) runtime_bd;
} MirrorRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(35)) matchtable_read_mirror(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_mirror(Bit#(18) msgtype, Bit#(35) data);
`endif
instance MatchTableSim#(104, 18, 35);
  function ActionValue#(Bit#(35)) matchtable_read(Bit#(104) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_mirror(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(104) id, Bit#(18) key, Bit#(35) data);
    action
      matchtable_write_mirror(key, data);
    endaction
  endfunction

endinstance
interface Mirror;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
endinterface
(* synthesize *)
module mkMirror  (Mirror);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(4, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(4, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(104, 1024, SizeOf#(MirrorReqT), SizeOf#(MirrorRspT)) matchTable <- mkMatchTable("mirror.dat");
  Vector#(4, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(4) readyChannel = -1;
  for (Integer i=3; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i2e_metadata$mirror_session_id = fromMaybe(?, meta.i2e_metadata$mirror_session_id);
    MirrorReqT req = MirrorReqT {i2e_metadata$mirror_session_id: i2e_metadata$mirror_session_id};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      MirrorRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_MIRROR_NHOP: begin
          BBRequest req = tagged SetMirrorNhopReqT {pkt: pkt, runtime_nhop_idx: resp.runtime_nhop_idx};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_MIRROR_BD: begin
          BBRequest req = tagged SetMirrorBdReqT {pkt: pkt, runtime_bd: resp.runtime_bd};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        SFLOW_PKT_TO_CPU: begin
          BBRequest req = tagged SflowPktToCpuReqT {pkt: pkt, sflow_metadata$sflow_session_id: sflow_metadata$sflow_session_id};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged MirrorNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMirrorNhopRspT {pkt: .pkt, l3_metadata$nexthop_index: .l3_metadata$nexthop_index}: begin
        meta.l3_metadata$nexthop_index = tagged Valid l3_metadata$nexthop_index;
        MetadataResponse rsp = tagged MirrorSetMirrorNhopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMirrorBdRspT {pkt: .pkt, egress_metadata$bd: .egress_metadata$bd}: begin
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        MetadataResponse rsp = tagged MirrorSetMirrorBdRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SflowPktToCpuRspT {pkt: .pkt, fabric_header_sflow$sflow_session_id: .fabric_header_sflow$sflow_session_id}: begin
        meta.fabric_header_sflow$sflow_session_id = tagged Valid fabric_header_sflow$sflow_session_id;
        MetadataResponse rsp = tagged MirrorSflowPktToCpuRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
endmodule

// ====== MTU ======

typedef struct {
  Bit#(8) padding;
  Bit#(8) l3_metadata$mtu_index;
  Bit#(Bool) valid_ipv4;
  Bit#(Bool) valid_ipv6;
} MtuReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_MTU,
  MTU_MISS,
  IPV4_MTU_CHECK,
  IPV6_MTU_CHECK
} MtuActionT deriving (Bits, Eq, FShow);
typedef struct {
  MtuActionT _action;
  Bit#(16) runtime_l3_mtu;
} MtuRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_mtu(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_mtu(Bit#(18) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(85, 18, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(85) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_mtu(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(85) id, Bit#(18) key, Bit#(18) data);
    action
      matchtable_write_mtu(key, data);
    endaction
  endfunction

endinstance
interface Mtu;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkMtu  (Mtu);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(85, 1024, SizeOf#(MtuReqT), SizeOf#(MtuRspT)) matchTable <- mkMatchTable("mtu.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$mtu_index = fromMaybe(?, meta.l3_metadata$mtu_index);
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let i$p$v$6 = fromMaybe(?, meta.i$p$v$6);
    MtuReqT req = MtuReqT {l3_metadata$mtu_index: l3_metadata$mtu_index,i$p$v$4: i$p$v$4,i$p$v$6: i$p$v$6};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      MtuRspT resp = unpack(data);
      case (resp._action) matches
        MTU_MISS: begin
          BBRequest req = tagged MtuMissReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_MTU_CHECK: begin
          BBRequest req = tagged Ipv4MtuCheckReqT {pkt: pkt, runtime_l3_mtu: resp.runtime_l3_mtu};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_MTU_CHECK: begin
          BBRequest req = tagged Ipv6MtuCheckReqT {pkt: pkt, runtime_l3_mtu: resp.runtime_l3_mtu};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged MtuMissRspT {pkt: .pkt, l3_metadata$l3_mtu_check: .l3_metadata$l3_mtu_check}: begin
        meta.l3_metadata$l3_mtu_check = tagged Valid l3_metadata$l3_mtu_check;
        MetadataResponse rsp = tagged MtuMtuMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4MtuCheckRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged MtuIpv4MtuCheckRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6MtuCheckRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged MtuIpv6MtuCheckRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== REPLICA_TYPE ======

typedef struct {
  Bit#(1) padding;
  Bit#(1) multicast_metadata$replica;
  Bit#(16) egress_metadata$same_bd_check;
} ReplicaTypeReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_REPLICA_TYPE,
  NOP,
  SET_REPLICA_COPY_BRIDGED
} ReplicaTypeActionT deriving (Bits, Eq, FShow);
typedef struct {
  ReplicaTypeActionT _action;
} ReplicaTypeRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_replica_type(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_replica_type(Bit#(18) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(99, 18, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(99) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_replica_type(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(99) id, Bit#(18) key, Bit#(2) data);
    action
      matchtable_write_replica_type(key, data);
    endaction
  endfunction

endinstance
interface ReplicaType;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkReplicaType  (ReplicaType);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(99, 512, SizeOf#(ReplicaTypeReqT), SizeOf#(ReplicaTypeRspT)) matchTable <- mkMatchTable("replica_type.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let multicast_metadata$replica = fromMaybe(?, meta.multicast_metadata$replica);
    let egress_metadata$same_bd_check = fromMaybe(?, meta.egress_metadata$same_bd_check);
    ReplicaTypeReqT req = ReplicaTypeReqT {multicast_metadata$replica: multicast_metadata$replica,egress_metadata$same_bd_check: egress_metadata$same_bd_check};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      ReplicaTypeRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_REPLICA_COPY_BRIDGED: begin
          BBRequest req = tagged SetReplicaCopyBridgedReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged ReplicaTypeNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetReplicaCopyBridgedRspT {pkt: .pkt, egress_metadata$routed: .egress_metadata$routed}: begin
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        MetadataResponse rsp = tagged ReplicaTypeSetReplicaCopyBridgedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== REWRITE ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) l3_metadata$nexthop_index;
} RewriteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_REWRITE,
  NOP,
  SET_L2_REWRITE,
  SET_L2_REWRITE_WITH_TUNNEL,
  SET_L3_REWRITE,
  SET_L3_REWRITE_WITH_TUNNEL,
  SET_MPLS_SWAP_PUSH_REWRITE_L2,
  SET_MPLS_PUSH_REWRITE_L2,
  SET_MPLS_SWAP_PUSH_REWRITE_L3,
  SET_MPLS_PUSH_REWRITE_L3
} RewriteActionT deriving (Bits, Eq, FShow);
typedef struct {
  RewriteActionT _action;
  Bit#(14) runtime_tunnel_index;
  Bit#(5) runtime_tunnel_type;
  Bit#(16) runtime_bd;
  Bit#(8) runtime_mtu_index;
  Bit#(48) runtime_dmac;
  Bit#(20) runtime_label;
  Bit#(4) runtime_header_count;
} RewriteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(119)) matchtable_read_rewrite(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_rewrite(Bit#(18) msgtype, Bit#(119) data);
`endif
instance MatchTableSim#(100, 18, 119);
  function ActionValue#(Bit#(119)) matchtable_read(Bit#(100) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_rewrite(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(100) id, Bit#(18) key, Bit#(119) data);
    action
      matchtable_write_rewrite(key, data);
    endaction
  endfunction

endinstance
interface Rewrite;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
endinterface
(* synthesize *)
module mkRewrite  (Rewrite);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(9, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(9, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(100, 1024, SizeOf#(RewriteReqT), SizeOf#(RewriteRspT)) matchTable <- mkMatchTable("rewrite.dat");
  Vector#(9, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(9) readyChannel = -1;
  for (Integer i=8; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
    RewriteReqT req = RewriteReqT {l3_metadata$nexthop_index: l3_metadata$nexthop_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      RewriteRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_L2_REWRITE: begin
          BBRequest req = tagged SetL2RewriteReqT {pkt: pkt, ingress_metadata$bd: ingress_metadata$bd};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_L2_REWRITE_WITH_TUNNEL: begin
          BBRequest req = tagged SetL2RewriteWithTunnelReqT {pkt: pkt, ingress_metadata$bd: ingress_metadata$bd, runtime_tunnel_index: resp.runtime_tunnel_index, runtime_tunnel_type: resp.runtime_tunnel_type};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        SET_L3_REWRITE: begin
          BBRequest req = tagged SetL3RewriteReqT {pkt: pkt, runtime_dmac: resp.runtime_dmac, runtime_bd: resp.runtime_bd, runtime_mtu_index: resp.runtime_mtu_index};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        SET_L3_REWRITE_WITH_TUNNEL: begin
          BBRequest req = tagged SetL3RewriteWithTunnelReqT {pkt: pkt, runtime_dmac: resp.runtime_dmac, runtime_tunnel_index: resp.runtime_tunnel_index, runtime_bd: resp.runtime_bd, runtime_tunnel_type: resp.runtime_tunnel_type};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        SET_MPLS_SWAP_PUSH_REWRITE_L2: begin
          BBRequest req = tagged SetMplsSwapPushRewriteL2ReqT {pkt: pkt, l3_metadata$routed: l3_metadata$routed, ingress_metadata$bd: ingress_metadata$bd, runtime_tunnel_index: resp.runtime_tunnel_index, runtime_label: resp.runtime_label, runtime_header_count: resp.runtime_header_count};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        SET_MPLS_PUSH_REWRITE_L2: begin
          BBRequest req = tagged SetMplsPushRewriteL2ReqT {pkt: pkt, l3_metadata$routed: l3_metadata$routed, ingress_metadata$bd: ingress_metadata$bd, runtime_tunnel_index: resp.runtime_tunnel_index, runtime_header_count: resp.runtime_header_count};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        SET_MPLS_SWAP_PUSH_REWRITE_L3: begin
          BBRequest req = tagged SetMplsSwapPushRewriteL3ReqT {pkt: pkt, l3_metadata$routed: l3_metadata$routed, runtime_dmac: resp.runtime_dmac, runtime_tunnel_index: resp.runtime_tunnel_index, runtime_label: resp.runtime_label, runtime_bd: resp.runtime_bd, runtime_header_count: resp.runtime_header_count};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        SET_MPLS_PUSH_REWRITE_L3: begin
          BBRequest req = tagged SetMplsPushRewriteL3ReqT {pkt: pkt, l3_metadata$routed: l3_metadata$routed, runtime_dmac: resp.runtime_dmac, runtime_tunnel_index: resp.runtime_tunnel_index, runtime_bd: resp.runtime_bd, runtime_header_count: resp.runtime_header_count};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged RewriteNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetL2RewriteRspT {pkt: .pkt, egress_metadata$outer_bd: .egress_metadata$outer_bd, egress_metadata$bd: .egress_metadata$bd, egress_metadata$routed: .egress_metadata$routed}: begin
        meta.egress_metadata$outer_bd = tagged Valid egress_metadata$outer_bd;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        MetadataResponse rsp = tagged RewriteSetL2RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetL2RewriteWithTunnelRspT {pkt: .pkt, egress_metadata$outer_bd: .egress_metadata$outer_bd, egress_metadata$bd: .egress_metadata$bd, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index, egress_metadata$routed: .egress_metadata$routed, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type}: begin
        meta.egress_metadata$outer_bd = tagged Valid egress_metadata$outer_bd;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        MetadataResponse rsp = tagged RewriteSetL2RewriteWithTunnelRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetL3RewriteRspT {pkt: .pkt, egress_metadata$outer_bd: .egress_metadata$outer_bd, egress_metadata$bd: .egress_metadata$bd, egress_metadata$mac_da: .egress_metadata$mac_da, egress_metadata$routed: .egress_metadata$routed, l3_metadata$mtu_index: .l3_metadata$mtu_index}: begin
        meta.egress_metadata$outer_bd = tagged Valid egress_metadata$outer_bd;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.egress_metadata$mac_da = tagged Valid egress_metadata$mac_da;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        meta.l3_metadata$mtu_index = tagged Valid l3_metadata$mtu_index;
        MetadataResponse rsp = tagged RewriteSetL3RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetL3RewriteWithTunnelRspT {pkt: .pkt, egress_metadata$outer_bd: .egress_metadata$outer_bd, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index, egress_metadata$mac_da: .egress_metadata$mac_da, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type, egress_metadata$bd: .egress_metadata$bd, egress_metadata$routed: .egress_metadata$routed}: begin
        meta.egress_metadata$outer_bd = tagged Valid egress_metadata$outer_bd;
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        meta.egress_metadata$mac_da = tagged Valid egress_metadata$mac_da;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        MetadataResponse rsp = tagged RewriteSetL3RewriteWithTunnelRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMplsSwapPushRewriteL2RspT {pkt: .pkt, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index, egress_metadata$routed: .egress_metadata$routed, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type, egress_metadata$bd: .egress_metadata$bd, tunnel_metadata$egress_header_count: .tunnel_metadata$egress_header_count, mpls0$label: .mpls0$label}: begin
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.tunnel_metadata$egress_header_count = tagged Valid tunnel_metadata$egress_header_count;
        meta.mpls0$label = tagged Valid mpls0$label;
        MetadataResponse rsp = tagged RewriteSetMplsSwapPushRewriteL2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMplsPushRewriteL2RspT {pkt: .pkt, egress_metadata$bd: .egress_metadata$bd, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index, tunnel_metadata$egress_header_count: .tunnel_metadata$egress_header_count, egress_metadata$routed: .egress_metadata$routed, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type}: begin
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        meta.tunnel_metadata$egress_header_count = tagged Valid tunnel_metadata$egress_header_count;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        MetadataResponse rsp = tagged RewriteSetMplsPushRewriteL2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMplsSwapPushRewriteL3RspT {pkt: .pkt, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index, tunnel_metadata$egress_header_count: .tunnel_metadata$egress_header_count, egress_metadata$mac_da: .egress_metadata$mac_da, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type, egress_metadata$bd: .egress_metadata$bd, egress_metadata$routed: .egress_metadata$routed, mpls0$label: .mpls0$label}: begin
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        meta.tunnel_metadata$egress_header_count = tagged Valid tunnel_metadata$egress_header_count;
        meta.egress_metadata$mac_da = tagged Valid egress_metadata$mac_da;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        meta.mpls0$label = tagged Valid mpls0$label;
        MetadataResponse rsp = tagged RewriteSetMplsSwapPushRewriteL3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMplsPushRewriteL3RspT {pkt: .pkt, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index, egress_metadata$routed: .egress_metadata$routed, egress_metadata$mac_da: .egress_metadata$mac_da, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type, egress_metadata$bd: .egress_metadata$bd, tunnel_metadata$egress_header_count: .tunnel_metadata$egress_header_count}: begin
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        meta.egress_metadata$mac_da = tagged Valid egress_metadata$mac_da;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.tunnel_metadata$egress_header_count = tagged Valid tunnel_metadata$egress_header_count;
        MetadataResponse rsp = tagged RewriteSetMplsPushRewriteL3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
endmodule

// ====== REWRITE_MULTICAST ======

typedef struct {
  Bit#(Bool) valid_ipv4;
  Bit#(Bool) valid_ipv6;
  Bit#(32) ipv4$dstAddr;
  Bit#(128) ipv6$dstAddr;
} RewriteMulticastReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_REWRITE_MULTICAST,
  NOP,
  REWRITE_IPV4_MULTICAST,
  REWRITE_IPV6_MULTICAST
} RewriteMulticastActionT deriving (Bits, Eq, FShow);
typedef struct {
  RewriteMulticastActionT _action;
} RewriteMulticastRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_rewrite_multicast(Bit#(162) msgtype);
import "BDPI" function Action matchtable_write_rewrite_multicast(Bit#(162) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(101, 162, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(101) id, Bit#(162) key);
    actionvalue
      let v <- matchtable_read_rewrite_multicast(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(101) id, Bit#(162) key, Bit#(2) data);
    action
      matchtable_write_rewrite_multicast(key, data);
    endaction
  endfunction

endinstance
interface RewriteMulticast;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkRewriteMulticast  (RewriteMulticast);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(101, 256, SizeOf#(RewriteMulticastReqT), SizeOf#(RewriteMulticastRspT)) matchTable <- mkMatchTable("rewrite_multicast.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let i$p$v$6 = fromMaybe(?, meta.i$p$v$6);
    let ipv4$dstAddr = fromMaybe(?, meta.ipv4$dstAddr);
    let ipv6$dstAddr = fromMaybe(?, meta.ipv6$dstAddr);
    RewriteMulticastReqT req = RewriteMulticastReqT {i$p$v$4: i$p$v$4,i$p$v$6: i$p$v$6,ipv4$dstAddr: ipv4$dstAddr,ipv6$dstAddr: ipv6$dstAddr};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      RewriteMulticastRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        REWRITE_IPV4_MULTICAST: begin
          BBRequest req = tagged RewriteIpv4MulticastReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        REWRITE_IPV6_MULTICAST: begin
          BBRequest req = tagged RewriteIpv6MulticastReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged RewriteMulticastNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RewriteIpv4MulticastRspT {pkt: .pkt, ethernet$dstAddr: .ethernet$dstAddr}: begin
        meta.ethernet$dstAddr = tagged Valid ethernet$dstAddr;
        MetadataResponse rsp = tagged RewriteMulticastRewriteIpv4MulticastRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RewriteIpv6MulticastRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged RewriteMulticastRewriteIpv6MulticastRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== RID ======

typedef struct {
  Bit#(2) padding;
  Bit#(16) intrinsic_metadata$egress_rid;
} RidReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_RID,
  NOP,
  OUTER_REPLICA_FROM_RID,
  INNER_REPLICA_FROM_RID
} RidActionT deriving (Bits, Eq, FShow);
typedef struct {
  RidActionT _action;
  Bit#(16) runtime_bd;
  Bit#(14) runtime_tunnel_index;
  Bit#(5) runtime_tunnel_type;
  Bit#(4) runtime_header_count;
} RidRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(41)) matchtable_read_rid(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_rid(Bit#(18) msgtype, Bit#(41) data);
`endif
instance MatchTableSim#(98, 18, 41);
  function ActionValue#(Bit#(41)) matchtable_read(Bit#(98) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_rid(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(98) id, Bit#(18) key, Bit#(41) data);
    action
      matchtable_write_rid(key, data);
    endaction
  endfunction

endinstance
interface Rid;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkRid  (Rid);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(98, 1024, SizeOf#(RidReqT), SizeOf#(RidRspT)) matchTable <- mkMatchTable("rid.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let intrinsic_metadata$egress_rid = fromMaybe(?, meta.intrinsic_metadata$egress_rid);
    RidReqT req = RidReqT {intrinsic_metadata$egress_rid: intrinsic_metadata$egress_rid};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      RidRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        OUTER_REPLICA_FROM_RID: begin
          BBRequest req = tagged OuterReplicaFromRidReqT {pkt: pkt, l3_metadata$outer_routed: l3_metadata$outer_routed, runtime_tunnel_index: resp.runtime_tunnel_index, runtime_tunnel_type: resp.runtime_tunnel_type, runtime_bd: resp.runtime_bd, runtime_header_count: resp.runtime_header_count};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        INNER_REPLICA_FROM_RID: begin
          BBRequest req = tagged InnerReplicaFromRidReqT {pkt: pkt, l3_metadata$routed: l3_metadata$routed, runtime_tunnel_index: resp.runtime_tunnel_index, runtime_tunnel_type: resp.runtime_tunnel_type, runtime_bd: resp.runtime_bd, runtime_header_count: resp.runtime_header_count};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged RidNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged OuterReplicaFromRidRspT {pkt: .pkt, multicast_metadata$replica: .multicast_metadata$replica, multicast_metadata$inner_replica: .multicast_metadata$inner_replica, tunnel_metadata$egress_header_count: .tunnel_metadata$egress_header_count, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type, egress_metadata$bd: .egress_metadata$bd, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index, egress_metadata$routed: .egress_metadata$routed}: begin
        meta.multicast_metadata$replica = tagged Valid multicast_metadata$replica;
        meta.multicast_metadata$inner_replica = tagged Valid multicast_metadata$inner_replica;
        meta.tunnel_metadata$egress_header_count = tagged Valid tunnel_metadata$egress_header_count;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        MetadataResponse rsp = tagged RidOuterReplicaFromRidRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerReplicaFromRidRspT {pkt: .pkt, multicast_metadata$replica: .multicast_metadata$replica, multicast_metadata$inner_replica: .multicast_metadata$inner_replica, tunnel_metadata$egress_header_count: .tunnel_metadata$egress_header_count, tunnel_metadata$egress_tunnel_type: .tunnel_metadata$egress_tunnel_type, egress_metadata$bd: .egress_metadata$bd, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index, egress_metadata$routed: .egress_metadata$routed}: begin
        meta.multicast_metadata$replica = tagged Valid multicast_metadata$replica;
        meta.multicast_metadata$inner_replica = tagged Valid multicast_metadata$inner_replica;
        meta.tunnel_metadata$egress_header_count = tagged Valid tunnel_metadata$egress_header_count;
        meta.tunnel_metadata$egress_tunnel_type = tagged Valid tunnel_metadata$egress_tunnel_type;
        meta.egress_metadata$bd = tagged Valid egress_metadata$bd;
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        meta.egress_metadata$routed = tagged Valid egress_metadata$routed;
        MetadataResponse rsp = tagged RidInnerReplicaFromRidRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== SMAC_REWRITE ======

typedef struct {
  Bit#(9) egress_metadata$smac_idx;
} SmacRewriteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_SMAC_REWRITE,
  REWRITE_SMAC
} SmacRewriteActionT deriving (Bits, Eq, FShow);
typedef struct {
  SmacRewriteActionT _action;
  Bit#(48) runtime_smac;
} SmacRewriteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(49)) matchtable_read_smac_rewrite(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_smac_rewrite(Bit#(9) msgtype, Bit#(49) data);
`endif
instance MatchTableSim#(83, 9, 49);
  function ActionValue#(Bit#(49)) matchtable_read(Bit#(83) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_smac_rewrite(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(83) id, Bit#(9) key, Bit#(49) data);
    action
      matchtable_write_smac_rewrite(key, data);
    endaction
  endfunction

endinstance
interface SmacRewrite;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
endinterface
(* synthesize *)
module mkSmacRewrite  (SmacRewrite);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(1, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(1, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(83, 512, SizeOf#(SmacRewriteReqT), SizeOf#(SmacRewriteRspT)) matchTable <- mkMatchTable("smac_rewrite.dat");
  Vector#(1, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(1) readyChannel = -1;
  for (Integer i=0; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let egress_metadata$smac_idx = fromMaybe(?, meta.egress_metadata$smac_idx);
    SmacRewriteReqT req = SmacRewriteReqT {egress_metadata$smac_idx: egress_metadata$smac_idx};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      SmacRewriteRspT resp = unpack(data);
      case (resp._action) matches
        REWRITE_SMAC: begin
          BBRequest req = tagged RewriteSmacReqT {pkt: pkt, runtime_smac: resp.runtime_smac};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged RewriteSmacRspT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr}: begin
        meta.ethernet$srcAddr = tagged Valid ethernet$srcAddr;
        MetadataResponse rsp = tagged SmacRewriteRewriteSmacRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
endmodule

// ====== TUNNEL_DECAP_PROCESS_INNER ======

typedef struct {
  Bit#(6) padding;
  Bit#(Bool) valid_inner_tcp;
  Bit#(Bool) valid_inner_udp;
  Bit#(Bool) valid_inner_icmp;
} TunnelDecapProcessInnerReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_DECAP_PROCESS_INNER,
  DECAP_INNER_UDP,
  DECAP_INNER_TCP,
  DECAP_INNER_ICMP,
  DECAP_INNER_UNKNOWN
} TunnelDecapProcessInnerActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelDecapProcessInnerActionT _action;
} TunnelDecapProcessInnerRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(3)) matchtable_read_tunnel_decap_process_inner(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_tunnel_decap_process_inner(Bit#(9) msgtype, Bit#(3) data);
`endif
instance MatchTableSim#(87, 9, 3);
  function ActionValue#(Bit#(3)) matchtable_read(Bit#(87) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_tunnel_decap_process_inner(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(87) id, Bit#(9) key, Bit#(3) data);
    action
      matchtable_write_tunnel_decap_process_inner(key, data);
    endaction
  endfunction

endinstance
interface TunnelDecapProcessInner;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
endinterface
(* synthesize *)
module mkTunnelDecapProcessInner  (TunnelDecapProcessInner);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(4, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(4, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(87, 1024, SizeOf#(TunnelDecapProcessInnerReqT), SizeOf#(TunnelDecapProcessInnerRspT)) matchTable <- mkMatchTable("tunnel_decap_process_inner.dat");
  Vector#(4, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(4) readyChannel = -1;
  for (Integer i=3; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$n$n$e$r$_$t$c$p = fromMaybe(?, meta.i$n$n$e$r$_$t$c$p);
    let i$n$n$e$r$_$u$d$p = fromMaybe(?, meta.i$n$n$e$r$_$u$d$p);
    let i$n$n$e$r$_$i$c$m$p = fromMaybe(?, meta.i$n$n$e$r$_$i$c$m$p);
    TunnelDecapProcessInnerReqT req = TunnelDecapProcessInnerReqT {i$n$n$e$r$_$t$c$p: i$n$n$e$r$_$t$c$p,i$n$n$e$r$_$u$d$p: i$n$n$e$r$_$u$d$p,i$n$n$e$r$_$i$c$m$p: i$n$n$e$r$_$i$c$m$p};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelDecapProcessInnerRspT resp = unpack(data);
      case (resp._action) matches
        DECAP_INNER_UDP: begin
          BBRequest req = tagged DecapInnerUdpReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_INNER_TCP: begin
          BBRequest req = tagged DecapInnerTcpReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_INNER_ICMP: begin
          BBRequest req = tagged DecapInnerIcmpReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_INNER_UNKNOWN: begin
          BBRequest req = tagged DecapInnerUnknownReqT {pkt: pkt};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged DecapInnerUdpRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessInnerDecapInnerUdpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapInnerTcpRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessInnerDecapInnerTcpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapInnerIcmpRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessInnerDecapInnerIcmpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapInnerUnknownRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessInnerDecapInnerUnknownRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
endmodule

// ====== TUNNEL_DECAP_PROCESS_OUTER ======

typedef struct {
  Bit#(2) padding;
  Bit#(5) tunnel_metadata$ingress_tunnel_type;
  Bit#(Bool) valid_inner_ipv4;
  Bit#(Bool) valid_inner_ipv6;
} TunnelDecapProcessOuterReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_DECAP_PROCESS_OUTER,
  DECAP_VXLAN_INNER_IPV4,
  DECAP_VXLAN_INNER_IPV6,
  DECAP_VXLAN_INNER_NON_IP,
  DECAP_GENV_INNER_IPV4,
  DECAP_GENV_INNER_IPV6,
  DECAP_GENV_INNER_NON_IP,
  DECAP_NVGRE_INNER_IPV4,
  DECAP_NVGRE_INNER_IPV6,
  DECAP_NVGRE_INNER_NON_IP,
  DECAP_GRE_INNER_IPV4,
  DECAP_GRE_INNER_IPV6,
  DECAP_GRE_INNER_NON_IP,
  DECAP_IP_INNER_IPV4,
  DECAP_IP_INNER_IPV6,
  DECAP_MPLS_INNER_IPV4_POP1,
  DECAP_MPLS_INNER_IPV6_POP1,
  DECAP_MPLS_INNER_ETHERNET_IPV4_POP1,
  DECAP_MPLS_INNER_ETHERNET_IPV6_POP1,
  DECAP_MPLS_INNER_ETHERNET_NON_IP_POP1,
  DECAP_MPLS_INNER_IPV4_POP2,
  DECAP_MPLS_INNER_IPV6_POP2,
  DECAP_MPLS_INNER_ETHERNET_IPV4_POP2,
  DECAP_MPLS_INNER_ETHERNET_IPV6_POP2,
  DECAP_MPLS_INNER_ETHERNET_NON_IP_POP2,
  DECAP_MPLS_INNER_IPV4_POP3,
  DECAP_MPLS_INNER_IPV6_POP3,
  DECAP_MPLS_INNER_ETHERNET_IPV4_POP3,
  DECAP_MPLS_INNER_ETHERNET_IPV6_POP3,
  DECAP_MPLS_INNER_ETHERNET_NON_IP_POP3
} TunnelDecapProcessOuterActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelDecapProcessOuterActionT _action;
} TunnelDecapProcessOuterRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(5)) matchtable_read_tunnel_decap_process_outer(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_tunnel_decap_process_outer(Bit#(9) msgtype, Bit#(5) data);
`endif
instance MatchTableSim#(86, 9, 5);
  function ActionValue#(Bit#(5)) matchtable_read(Bit#(86) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_tunnel_decap_process_outer(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(86) id, Bit#(9) key, Bit#(5) data);
    action
      matchtable_write_tunnel_decap_process_outer(key, data);
    endaction
  endfunction

endinstance
interface TunnelDecapProcessOuter;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
  interface Client #(BBRequest, BBResponse) next_control_state_9;
  interface Client #(BBRequest, BBResponse) next_control_state_10;
  interface Client #(BBRequest, BBResponse) next_control_state_11;
  interface Client #(BBRequest, BBResponse) next_control_state_12;
  interface Client #(BBRequest, BBResponse) next_control_state_13;
  interface Client #(BBRequest, BBResponse) next_control_state_14;
  interface Client #(BBRequest, BBResponse) next_control_state_15;
  interface Client #(BBRequest, BBResponse) next_control_state_16;
  interface Client #(BBRequest, BBResponse) next_control_state_17;
  interface Client #(BBRequest, BBResponse) next_control_state_18;
  interface Client #(BBRequest, BBResponse) next_control_state_19;
  interface Client #(BBRequest, BBResponse) next_control_state_20;
  interface Client #(BBRequest, BBResponse) next_control_state_21;
  interface Client #(BBRequest, BBResponse) next_control_state_22;
  interface Client #(BBRequest, BBResponse) next_control_state_23;
  interface Client #(BBRequest, BBResponse) next_control_state_24;
  interface Client #(BBRequest, BBResponse) next_control_state_25;
  interface Client #(BBRequest, BBResponse) next_control_state_26;
  interface Client #(BBRequest, BBResponse) next_control_state_27;
  interface Client #(BBRequest, BBResponse) next_control_state_28;
endinterface
(* synthesize *)
module mkTunnelDecapProcessOuter  (TunnelDecapProcessOuter);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(29, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(29, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(86, 1024, SizeOf#(TunnelDecapProcessOuterReqT), SizeOf#(TunnelDecapProcessOuterRspT)) matchTable <- mkMatchTable("tunnel_decap_process_outer.dat");
  Vector#(29, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(29) readyChannel = -1;
  for (Integer i=28; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
    let i$n$n$e$r$_$i$p$v$4 = fromMaybe(?, meta.i$n$n$e$r$_$i$p$v$4);
    let i$n$n$e$r$_$i$p$v$6 = fromMaybe(?, meta.i$n$n$e$r$_$i$p$v$6);
    TunnelDecapProcessOuterReqT req = TunnelDecapProcessOuterReqT {tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type,i$n$n$e$r$_$i$p$v$4: i$n$n$e$r$_$i$p$v$4,i$n$n$e$r$_$i$p$v$6: i$n$n$e$r$_$i$p$v$6};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelDecapProcessOuterRspT resp = unpack(data);
      case (resp._action) matches
        DECAP_VXLAN_INNER_IPV4: begin
          BBRequest req = tagged DecapVxlanInnerIpv4ReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_VXLAN_INNER_IPV6: begin
          BBRequest req = tagged DecapVxlanInnerIpv6ReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_VXLAN_INNER_NON_IP: begin
          BBRequest req = tagged DecapVxlanInnerNonIpReqT {pkt: pkt};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_GENV_INNER_IPV4: begin
          BBRequest req = tagged DecapGenvInnerIpv4ReqT {pkt: pkt};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_GENV_INNER_IPV6: begin
          BBRequest req = tagged DecapGenvInnerIpv6ReqT {pkt: pkt};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_GENV_INNER_NON_IP: begin
          BBRequest req = tagged DecapGenvInnerNonIpReqT {pkt: pkt};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_NVGRE_INNER_IPV4: begin
          BBRequest req = tagged DecapNvgreInnerIpv4ReqT {pkt: pkt};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_NVGRE_INNER_IPV6: begin
          BBRequest req = tagged DecapNvgreInnerIpv6ReqT {pkt: pkt};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_NVGRE_INNER_NON_IP: begin
          BBRequest req = tagged DecapNvgreInnerNonIpReqT {pkt: pkt};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_GRE_INNER_IPV4: begin
          BBRequest req = tagged DecapGreInnerIpv4ReqT {pkt: pkt};
          bbReqFifo[9].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_GRE_INNER_IPV6: begin
          BBRequest req = tagged DecapGreInnerIpv6ReqT {pkt: pkt};
          bbReqFifo[10].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_GRE_INNER_NON_IP: begin
          BBRequest req = tagged DecapGreInnerNonIpReqT {pkt: pkt, gre$proto: gre$proto};
          bbReqFifo[11].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_IP_INNER_IPV4: begin
          BBRequest req = tagged DecapIpInnerIpv4ReqT {pkt: pkt};
          bbReqFifo[12].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_IP_INNER_IPV6: begin
          BBRequest req = tagged DecapIpInnerIpv6ReqT {pkt: pkt};
          bbReqFifo[13].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_IPV4_POP1: begin
          BBRequest req = tagged DecapMplsInnerIpv4Pop1ReqT {pkt: pkt};
          bbReqFifo[14].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_IPV6_POP1: begin
          BBRequest req = tagged DecapMplsInnerIpv6Pop1ReqT {pkt: pkt};
          bbReqFifo[15].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_IPV4_POP1: begin
          BBRequest req = tagged DecapMplsInnerEthernetIpv4Pop1ReqT {pkt: pkt};
          bbReqFifo[16].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_IPV6_POP1: begin
          BBRequest req = tagged DecapMplsInnerEthernetIpv6Pop1ReqT {pkt: pkt};
          bbReqFifo[17].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_NON_IP_POP1: begin
          BBRequest req = tagged DecapMplsInnerEthernetNonIpPop1ReqT {pkt: pkt};
          bbReqFifo[18].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_IPV4_POP2: begin
          BBRequest req = tagged DecapMplsInnerIpv4Pop2ReqT {pkt: pkt};
          bbReqFifo[19].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_IPV6_POP2: begin
          BBRequest req = tagged DecapMplsInnerIpv6Pop2ReqT {pkt: pkt};
          bbReqFifo[20].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_IPV4_POP2: begin
          BBRequest req = tagged DecapMplsInnerEthernetIpv4Pop2ReqT {pkt: pkt};
          bbReqFifo[21].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_IPV6_POP2: begin
          BBRequest req = tagged DecapMplsInnerEthernetIpv6Pop2ReqT {pkt: pkt};
          bbReqFifo[22].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_NON_IP_POP2: begin
          BBRequest req = tagged DecapMplsInnerEthernetNonIpPop2ReqT {pkt: pkt};
          bbReqFifo[23].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_IPV4_POP3: begin
          BBRequest req = tagged DecapMplsInnerIpv4Pop3ReqT {pkt: pkt};
          bbReqFifo[24].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_IPV6_POP3: begin
          BBRequest req = tagged DecapMplsInnerIpv6Pop3ReqT {pkt: pkt};
          bbReqFifo[25].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_IPV4_POP3: begin
          BBRequest req = tagged DecapMplsInnerEthernetIpv4Pop3ReqT {pkt: pkt};
          bbReqFifo[26].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_IPV6_POP3: begin
          BBRequest req = tagged DecapMplsInnerEthernetIpv6Pop3ReqT {pkt: pkt};
          bbReqFifo[27].enq(req); //FIXME: replace with RXTX.
        end
        DECAP_MPLS_INNER_ETHERNET_NON_IP_POP3: begin
          BBRequest req = tagged DecapMplsInnerEthernetNonIpPop3ReqT {pkt: pkt};
          bbReqFifo[28].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged DecapVxlanInnerIpv4RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapVxlanInnerIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapVxlanInnerIpv6RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapVxlanInnerIpv6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapVxlanInnerNonIpRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapVxlanInnerNonIpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapGenvInnerIpv4RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapGenvInnerIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapGenvInnerIpv6RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapGenvInnerIpv6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapGenvInnerNonIpRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapGenvInnerNonIpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapNvgreInnerIpv4RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapNvgreInnerIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapNvgreInnerIpv6RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapNvgreInnerIpv6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapNvgreInnerNonIpRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapNvgreInnerNonIpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapGreInnerIpv4RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapGreInnerIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapGreInnerIpv6RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapGreInnerIpv6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapGreInnerNonIpRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapGreInnerNonIpRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapIpInnerIpv4RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapIpInnerIpv4RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapIpInnerIpv6RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapIpInnerIpv6RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerIpv4Pop1RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerIpv4Pop1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerIpv6Pop1RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerIpv6Pop1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetIpv4Pop1RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv4Pop1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetIpv6Pop1RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv6Pop1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetNonIpPop1RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetNonIpPop1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerIpv4Pop2RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerIpv4Pop2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerIpv6Pop2RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerIpv6Pop2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetIpv4Pop2RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv4Pop2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetIpv6Pop2RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv6Pop2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetNonIpPop2RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetNonIpPop2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerIpv4Pop3RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerIpv4Pop3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerIpv6Pop3RspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerIpv6Pop3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetIpv4Pop3RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv4Pop3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetIpv6Pop3RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv6Pop3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged DecapMplsInnerEthernetNonIpPop3RspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDecapProcessOuterDecapMplsInnerEthernetNonIpPop3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
  interface next_control_state_9 = toClient(bbReqFifo[9], bbRspFifo[9]);
  interface next_control_state_10 = toClient(bbReqFifo[10], bbRspFifo[10]);
  interface next_control_state_11 = toClient(bbReqFifo[11], bbRspFifo[11]);
  interface next_control_state_12 = toClient(bbReqFifo[12], bbRspFifo[12]);
  interface next_control_state_13 = toClient(bbReqFifo[13], bbRspFifo[13]);
  interface next_control_state_14 = toClient(bbReqFifo[14], bbRspFifo[14]);
  interface next_control_state_15 = toClient(bbReqFifo[15], bbRspFifo[15]);
  interface next_control_state_16 = toClient(bbReqFifo[16], bbRspFifo[16]);
  interface next_control_state_17 = toClient(bbReqFifo[17], bbRspFifo[17]);
  interface next_control_state_18 = toClient(bbReqFifo[18], bbRspFifo[18]);
  interface next_control_state_19 = toClient(bbReqFifo[19], bbRspFifo[19]);
  interface next_control_state_20 = toClient(bbReqFifo[20], bbRspFifo[20]);
  interface next_control_state_21 = toClient(bbReqFifo[21], bbRspFifo[21]);
  interface next_control_state_22 = toClient(bbReqFifo[22], bbRspFifo[22]);
  interface next_control_state_23 = toClient(bbReqFifo[23], bbRspFifo[23]);
  interface next_control_state_24 = toClient(bbReqFifo[24], bbRspFifo[24]);
  interface next_control_state_25 = toClient(bbReqFifo[25], bbRspFifo[25]);
  interface next_control_state_26 = toClient(bbReqFifo[26], bbRspFifo[26]);
  interface next_control_state_27 = toClient(bbReqFifo[27], bbRspFifo[27]);
  interface next_control_state_28 = toClient(bbReqFifo[28], bbRspFifo[28]);
endmodule

// ====== TUNNEL_DMAC_REWRITE ======

typedef struct {
  Bit#(4) padding;
  Bit#(14) tunnel_metadata$tunnel_dmac_index;
} TunnelDmacRewriteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_DMAC_REWRITE,
  NOP,
  REWRITE_TUNNEL_DMAC
} TunnelDmacRewriteActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelDmacRewriteActionT _action;
  Bit#(48) runtime_dmac;
} TunnelDmacRewriteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(50)) matchtable_read_tunnel_dmac_rewrite(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_tunnel_dmac_rewrite(Bit#(18) msgtype, Bit#(50) data);
`endif
instance MatchTableSim#(96, 18, 50);
  function ActionValue#(Bit#(50)) matchtable_read(Bit#(96) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_tunnel_dmac_rewrite(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(96) id, Bit#(18) key, Bit#(50) data);
    action
      matchtable_write_tunnel_dmac_rewrite(key, data);
    endaction
  endfunction

endinstance
interface TunnelDmacRewrite;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkTunnelDmacRewrite  (TunnelDmacRewrite);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(96, 1024, SizeOf#(TunnelDmacRewriteReqT), SizeOf#(TunnelDmacRewriteRspT)) matchTable <- mkMatchTable("tunnel_dmac_rewrite.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$tunnel_dmac_index = fromMaybe(?, meta.tunnel_metadata$tunnel_dmac_index);
    TunnelDmacRewriteReqT req = TunnelDmacRewriteReqT {tunnel_metadata$tunnel_dmac_index: tunnel_metadata$tunnel_dmac_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelDmacRewriteRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        REWRITE_TUNNEL_DMAC: begin
          BBRequest req = tagged RewriteTunnelDmacReqT {pkt: pkt, runtime_dmac: resp.runtime_dmac};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDmacRewriteNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RewriteTunnelDmacRspT {pkt: .pkt, ethernet$dstAddr: .ethernet$dstAddr}: begin
        meta.ethernet$dstAddr = tagged Valid ethernet$dstAddr;
        MetadataResponse rsp = tagged TunnelDmacRewriteRewriteTunnelDmacRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== TUNNEL_DST_REWRITE ======

typedef struct {
  Bit#(4) padding;
  Bit#(14) tunnel_metadata$tunnel_dst_index;
} TunnelDstRewriteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_DST_REWRITE,
  NOP,
  REWRITE_TUNNEL_IPV4_DST,
  REWRITE_TUNNEL_IPV6_DST
} TunnelDstRewriteActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelDstRewriteActionT _action;
  Bit#(32) runtime_ip;
} TunnelDstRewriteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_tunnel_dst_rewrite(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_tunnel_dst_rewrite(Bit#(18) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(94, 18, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(94) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_tunnel_dst_rewrite(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(94) id, Bit#(18) key, Bit#(34) data);
    action
      matchtable_write_tunnel_dst_rewrite(key, data);
    endaction
  endfunction

endinstance
interface TunnelDstRewrite;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkTunnelDstRewrite  (TunnelDstRewrite);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(94, 1024, SizeOf#(TunnelDstRewriteReqT), SizeOf#(TunnelDstRewriteRspT)) matchTable <- mkMatchTable("tunnel_dst_rewrite.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$tunnel_dst_index = fromMaybe(?, meta.tunnel_metadata$tunnel_dst_index);
    TunnelDstRewriteReqT req = TunnelDstRewriteReqT {tunnel_metadata$tunnel_dst_index: tunnel_metadata$tunnel_dst_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelDstRewriteRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        REWRITE_TUNNEL_IPV4_DST: begin
          BBRequest req = tagged RewriteTunnelIpv4DstReqT {pkt: pkt, runtime_ip: resp.runtime_ip};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        REWRITE_TUNNEL_IPV6_DST: begin
          BBRequest req = tagged RewriteTunnelIpv6DstReqT {pkt: pkt, runtime_ip: resp.runtime_ip};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelDstRewriteNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RewriteTunnelIpv4DstRspT {pkt: .pkt, ipv4$dstAddr: .ipv4$dstAddr}: begin
        meta.ipv4$dstAddr = tagged Valid ipv4$dstAddr;
        MetadataResponse rsp = tagged TunnelDstRewriteRewriteTunnelIpv4DstRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RewriteTunnelIpv6DstRspT {pkt: .pkt, ipv6$dstAddr: .ipv6$dstAddr}: begin
        meta.ipv6$dstAddr = tagged Valid ipv6$dstAddr;
        MetadataResponse rsp = tagged TunnelDstRewriteRewriteTunnelIpv6DstRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== TUNNEL_ENCAP_PROCESS_INNER ======

typedef struct {
  Bit#(4) padding;
  Bit#(Bool) valid_ipv4;
  Bit#(Bool) valid_ipv6;
  Bit#(Bool) valid_tcp;
  Bit#(Bool) valid_udp;
  Bit#(Bool) valid_icmp;
} TunnelEncapProcessInnerReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_ENCAP_PROCESS_INNER,
  INNER_IPV4_UDP_REWRITE,
  INNER_IPV4_TCP_REWRITE,
  INNER_IPV4_ICMP_REWRITE,
  INNER_IPV4_UNKNOWN_REWRITE,
  INNER_IPV6_UDP_REWRITE,
  INNER_IPV6_TCP_REWRITE,
  INNER_IPV6_ICMP_REWRITE,
  INNER_IPV6_UNKNOWN_REWRITE,
  INNER_NON_IP_REWRITE
} TunnelEncapProcessInnerActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelEncapProcessInnerActionT _action;
} TunnelEncapProcessInnerRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(4)) matchtable_read_tunnel_encap_process_inner(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_tunnel_encap_process_inner(Bit#(9) msgtype, Bit#(4) data);
`endif
instance MatchTableSim#(89, 9, 4);
  function ActionValue#(Bit#(4)) matchtable_read(Bit#(89) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_tunnel_encap_process_inner(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(89) id, Bit#(9) key, Bit#(4) data);
    action
      matchtable_write_tunnel_encap_process_inner(key, data);
    endaction
  endfunction

endinstance
interface TunnelEncapProcessInner;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
endinterface
(* synthesize *)
module mkTunnelEncapProcessInner  (TunnelEncapProcessInner);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(9, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(9, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(89, 1024, SizeOf#(TunnelEncapProcessInnerReqT), SizeOf#(TunnelEncapProcessInnerRspT)) matchTable <- mkMatchTable("tunnel_encap_process_inner.dat");
  Vector#(9, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(9) readyChannel = -1;
  for (Integer i=8; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let i$p$v$4 = fromMaybe(?, meta.i$p$v$4);
    let i$p$v$6 = fromMaybe(?, meta.i$p$v$6);
    let t$c$p = fromMaybe(?, meta.t$c$p);
    let u$d$p = fromMaybe(?, meta.u$d$p);
    let i$c$m$p = fromMaybe(?, meta.i$c$m$p);
    TunnelEncapProcessInnerReqT req = TunnelEncapProcessInnerReqT {i$p$v$4: i$p$v$4,i$p$v$6: i$p$v$6,t$c$p: t$c$p,u$d$p: u$d$p,i$c$m$p: i$c$m$p};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelEncapProcessInnerRspT resp = unpack(data);
      case (resp._action) matches
        INNER_IPV4_UDP_REWRITE: begin
          BBRequest req = tagged InnerIpv4UdpRewriteReqT {pkt: pkt, ipv4$totalLen: ipv4$totalLen};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        INNER_IPV4_TCP_REWRITE: begin
          BBRequest req = tagged InnerIpv4TcpRewriteReqT {pkt: pkt, ipv4$totalLen: ipv4$totalLen};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        INNER_IPV4_ICMP_REWRITE: begin
          BBRequest req = tagged InnerIpv4IcmpRewriteReqT {pkt: pkt, ipv4$totalLen: ipv4$totalLen};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        INNER_IPV4_UNKNOWN_REWRITE: begin
          BBRequest req = tagged InnerIpv4UnknownRewriteReqT {pkt: pkt, ipv4$totalLen: ipv4$totalLen};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        INNER_IPV6_UDP_REWRITE: begin
          BBRequest req = tagged InnerIpv6UdpRewriteReqT {pkt: pkt};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        INNER_IPV6_TCP_REWRITE: begin
          BBRequest req = tagged InnerIpv6TcpRewriteReqT {pkt: pkt};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        INNER_IPV6_ICMP_REWRITE: begin
          BBRequest req = tagged InnerIpv6IcmpRewriteReqT {pkt: pkt};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        INNER_IPV6_UNKNOWN_REWRITE: begin
          BBRequest req = tagged InnerIpv6UnknownRewriteReqT {pkt: pkt};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        INNER_NON_IP_REWRITE: begin
          BBRequest req = tagged InnerNonIpRewriteReqT {pkt: pkt};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged InnerIpv4UdpRewriteRspT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: .egress_metadata$payload_length}: begin
        meta.tunnel_metadata$inner_ip_proto = tagged Valid tunnel_metadata$inner_ip_proto;
        meta.egress_metadata$payload_length = tagged Valid egress_metadata$payload_length;
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerIpv4UdpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerIpv4TcpRewriteRspT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: .egress_metadata$payload_length}: begin
        meta.tunnel_metadata$inner_ip_proto = tagged Valid tunnel_metadata$inner_ip_proto;
        meta.egress_metadata$payload_length = tagged Valid egress_metadata$payload_length;
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerIpv4TcpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerIpv4IcmpRewriteRspT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: .egress_metadata$payload_length}: begin
        meta.tunnel_metadata$inner_ip_proto = tagged Valid tunnel_metadata$inner_ip_proto;
        meta.egress_metadata$payload_length = tagged Valid egress_metadata$payload_length;
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerIpv4IcmpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerIpv4UnknownRewriteRspT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: .egress_metadata$payload_length}: begin
        meta.tunnel_metadata$inner_ip_proto = tagged Valid tunnel_metadata$inner_ip_proto;
        meta.egress_metadata$payload_length = tagged Valid egress_metadata$payload_length;
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerIpv4UnknownRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerIpv6UdpRewriteRspT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto}: begin
        meta.tunnel_metadata$inner_ip_proto = tagged Valid tunnel_metadata$inner_ip_proto;
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerIpv6UdpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerIpv6TcpRewriteRspT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto}: begin
        meta.tunnel_metadata$inner_ip_proto = tagged Valid tunnel_metadata$inner_ip_proto;
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerIpv6TcpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerIpv6IcmpRewriteRspT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto}: begin
        meta.tunnel_metadata$inner_ip_proto = tagged Valid tunnel_metadata$inner_ip_proto;
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerIpv6IcmpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerIpv6UnknownRewriteRspT {pkt: .pkt, tunnel_metadata$inner_ip_proto: .tunnel_metadata$inner_ip_proto}: begin
        meta.tunnel_metadata$inner_ip_proto = tagged Valid tunnel_metadata$inner_ip_proto;
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerIpv6UnknownRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged InnerNonIpRewriteRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelEncapProcessInnerInnerNonIpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
endmodule

// ====== TUNNEL_ENCAP_PROCESS_OUTER ======

typedef struct {
  Bit#(8) padding;
  Bit#(5) tunnel_metadata$egress_tunnel_type;
  Bit#(4) tunnel_metadata$egress_header_count;
  Bit#(1) multicast_metadata$replica;
} TunnelEncapProcessOuterReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_ENCAP_PROCESS_OUTER,
  NOP,
  IPV4_VXLAN_REWRITE,
  IPV4_GENV_REWRITE,
  IPV4_NVGRE_REWRITE,
  IPV4_GRE_REWRITE,
  IPV4_IP_REWRITE,
  IPV4_ERSPAN_T3_REWRITE,
  IPV6_GRE_REWRITE,
  IPV6_IP_REWRITE,
  IPV6_NVGRE_REWRITE,
  IPV6_VXLAN_REWRITE,
  IPV6_GENV_REWRITE,
  IPV6_ERSPAN_T3_REWRITE,
  MPLS_ETHERNET_PUSH1_REWRITE,
  MPLS_IP_PUSH1_REWRITE,
  MPLS_ETHERNET_PUSH2_REWRITE,
  MPLS_IP_PUSH2_REWRITE,
  MPLS_ETHERNET_PUSH3_REWRITE,
  MPLS_IP_PUSH3_REWRITE,
  FABRIC_REWRITE
} TunnelEncapProcessOuterActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelEncapProcessOuterActionT _action;
  Bit#(14) runtime_tunnel_index;
} TunnelEncapProcessOuterRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(19)) matchtable_read_tunnel_encap_process_outer(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_tunnel_encap_process_outer(Bit#(18) msgtype, Bit#(19) data);
`endif
instance MatchTableSim#(90, 18, 19);
  function ActionValue#(Bit#(19)) matchtable_read(Bit#(90) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_tunnel_encap_process_outer(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(90) id, Bit#(18) key, Bit#(19) data);
    action
      matchtable_write_tunnel_encap_process_outer(key, data);
    endaction
  endfunction

endinstance
interface TunnelEncapProcessOuter;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
  interface Client #(BBRequest, BBResponse) next_control_state_8;
  interface Client #(BBRequest, BBResponse) next_control_state_9;
  interface Client #(BBRequest, BBResponse) next_control_state_10;
  interface Client #(BBRequest, BBResponse) next_control_state_11;
  interface Client #(BBRequest, BBResponse) next_control_state_12;
  interface Client #(BBRequest, BBResponse) next_control_state_13;
  interface Client #(BBRequest, BBResponse) next_control_state_14;
  interface Client #(BBRequest, BBResponse) next_control_state_15;
  interface Client #(BBRequest, BBResponse) next_control_state_16;
  interface Client #(BBRequest, BBResponse) next_control_state_17;
  interface Client #(BBRequest, BBResponse) next_control_state_18;
  interface Client #(BBRequest, BBResponse) next_control_state_19;
endinterface
(* synthesize *)
module mkTunnelEncapProcessOuter  (TunnelEncapProcessOuter);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(20, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(20, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(90, 1024, SizeOf#(TunnelEncapProcessOuterReqT), SizeOf#(TunnelEncapProcessOuterRspT)) matchTable <- mkMatchTable("tunnel_encap_process_outer.dat");
  Vector#(20, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(20) readyChannel = -1;
  for (Integer i=19; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
    let tunnel_metadata$egress_header_count = fromMaybe(?, meta.tunnel_metadata$egress_header_count);
    let multicast_metadata$replica = fromMaybe(?, meta.multicast_metadata$replica);
    TunnelEncapProcessOuterReqT req = TunnelEncapProcessOuterReqT {tunnel_metadata$egress_tunnel_type: tunnel_metadata$egress_tunnel_type,tunnel_metadata$egress_header_count: tunnel_metadata$egress_header_count,multicast_metadata$replica: multicast_metadata$replica};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelEncapProcessOuterRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_VXLAN_REWRITE: begin
          BBRequest req = tagged Ipv4VxlanRewriteReqT {pkt: pkt, hash_metadata$entropy_hash: hash_metadata$entropy_hash, tunnel_metadata$vnid: tunnel_metadata$vnid};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_GENV_REWRITE: begin
          BBRequest req = tagged Ipv4GenvRewriteReqT {pkt: pkt, hash_metadata$entropy_hash: hash_metadata$entropy_hash, tunnel_metadata$vnid: tunnel_metadata$vnid};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_NVGRE_REWRITE: begin
          BBRequest req = tagged Ipv4NvgreRewriteReqT {pkt: pkt, tunnel_metadata$vnid: tunnel_metadata$vnid};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_GRE_REWRITE: begin
          BBRequest req = tagged Ipv4GreRewriteReqT {pkt: pkt, ethernet$etherType: ethernet$etherType};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_IP_REWRITE: begin
          BBRequest req = tagged Ipv4IpRewriteReqT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        IPV4_ERSPAN_T3_REWRITE: begin
          BBRequest req = tagged Ipv4ErspanT3RewriteReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp, i2e_metadata$mirror_session_id: i2e_metadata$mirror_session_id};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_GRE_REWRITE: begin
          BBRequest req = tagged Ipv6GreRewriteReqT {pkt: pkt, ethernet$etherType: ethernet$etherType};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_IP_REWRITE: begin
          BBRequest req = tagged Ipv6IpRewriteReqT {pkt: pkt, tunnel_metadata$inner_ip_proto: tunnel_metadata$inner_ip_proto, egress_metadata$payload_length: egress_metadata$payload_length};
          bbReqFifo[8].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_NVGRE_REWRITE: begin
          BBRequest req = tagged Ipv6NvgreRewriteReqT {pkt: pkt, tunnel_metadata$vnid: tunnel_metadata$vnid};
          bbReqFifo[9].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_VXLAN_REWRITE: begin
          BBRequest req = tagged Ipv6VxlanRewriteReqT {pkt: pkt, hash_metadata$entropy_hash: hash_metadata$entropy_hash, tunnel_metadata$vnid: tunnel_metadata$vnid};
          bbReqFifo[10].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_GENV_REWRITE: begin
          BBRequest req = tagged Ipv6GenvRewriteReqT {pkt: pkt, hash_metadata$entropy_hash: hash_metadata$entropy_hash, tunnel_metadata$vnid: tunnel_metadata$vnid};
          bbReqFifo[11].enq(req); //FIXME: replace with RXTX.
        end
        IPV6_ERSPAN_T3_REWRITE: begin
          BBRequest req = tagged Ipv6ErspanT3RewriteReqT {pkt: pkt, i2e_metadata$ingress_tstamp: i2e_metadata$ingress_tstamp, i2e_metadata$mirror_session_id: i2e_metadata$mirror_session_id};
          bbReqFifo[12].enq(req); //FIXME: replace with RXTX.
        end
        MPLS_ETHERNET_PUSH1_REWRITE: begin
          BBRequest req = tagged MplsEthernetPush1RewriteReqT {pkt: pkt};
          bbReqFifo[13].enq(req); //FIXME: replace with RXTX.
        end
        MPLS_IP_PUSH1_REWRITE: begin
          BBRequest req = tagged MplsIpPush1RewriteReqT {pkt: pkt};
          bbReqFifo[14].enq(req); //FIXME: replace with RXTX.
        end
        MPLS_ETHERNET_PUSH2_REWRITE: begin
          BBRequest req = tagged MplsEthernetPush2RewriteReqT {pkt: pkt};
          bbReqFifo[15].enq(req); //FIXME: replace with RXTX.
        end
        MPLS_IP_PUSH2_REWRITE: begin
          BBRequest req = tagged MplsIpPush2RewriteReqT {pkt: pkt};
          bbReqFifo[16].enq(req); //FIXME: replace with RXTX.
        end
        MPLS_ETHERNET_PUSH3_REWRITE: begin
          BBRequest req = tagged MplsEthernetPush3RewriteReqT {pkt: pkt};
          bbReqFifo[17].enq(req); //FIXME: replace with RXTX.
        end
        MPLS_IP_PUSH3_REWRITE: begin
          BBRequest req = tagged MplsIpPush3RewriteReqT {pkt: pkt};
          bbReqFifo[18].enq(req); //FIXME: replace with RXTX.
        end
        FABRIC_REWRITE: begin
          BBRequest req = tagged FabricRewriteReqT {pkt: pkt, runtime_tunnel_index: resp.runtime_tunnel_index};
          bbReqFifo[19].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelEncapProcessOuterNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4VxlanRewriteRspT {pkt: .pkt, ipv4$identification: .ipv4$identification, udp$checksum: .udp$checksum, vxlan$vni: .vxlan$vni, ipv4$ihl: .ipv4$ihl, vxlan$flags: .vxlan$flags, ipv4$ttl: .ipv4$ttl, ipv4$protocol: .ipv4$protocol, vxlan$reserved2: .vxlan$reserved2, udp$srcPort: .udp$srcPort, vxlan$reserved: .vxlan$reserved, udp$dstPort: .udp$dstPort, ethernet$etherType: .ethernet$etherType, ipv4$version: .ipv4$version}: begin
        meta.ipv4$identification = tagged Valid ipv4$identification;
        meta.udp$checksum = tagged Valid udp$checksum;
        meta.vxlan$vni = tagged Valid vxlan$vni;
        meta.ipv4$ihl = tagged Valid ipv4$ihl;
        meta.vxlan$flags = tagged Valid vxlan$flags;
        meta.ipv4$ttl = tagged Valid ipv4$ttl;
        meta.ipv4$protocol = tagged Valid ipv4$protocol;
        meta.vxlan$reserved2 = tagged Valid vxlan$reserved2;
        meta.udp$srcPort = tagged Valid udp$srcPort;
        meta.vxlan$reserved = tagged Valid vxlan$reserved;
        meta.udp$dstPort = tagged Valid udp$dstPort;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.ipv4$version = tagged Valid ipv4$version;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv4VxlanRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4GenvRewriteRspT {pkt: .pkt, genv$vni: .genv$vni, ipv4$identification: .ipv4$identification, udp$checksum: .udp$checksum, ipv4$version: .ipv4$version, ipv4$ihl: .ipv4$ihl, genv$optLen: .genv$optLen, ipv4$ttl: .ipv4$ttl, genv$oam: .genv$oam, genv$reserved2: .genv$reserved2, genv$critical: .genv$critical, udp$srcPort: .udp$srcPort, genv$protoType: .genv$protoType, genv$ver: .genv$ver, udp$dstPort: .udp$dstPort, ethernet$etherType: .ethernet$etherType, ipv4$protocol: .ipv4$protocol, genv$reserved: .genv$reserved}: begin
        meta.genv$vni = tagged Valid genv$vni;
        meta.ipv4$identification = tagged Valid ipv4$identification;
        meta.udp$checksum = tagged Valid udp$checksum;
        meta.ipv4$version = tagged Valid ipv4$version;
        meta.ipv4$ihl = tagged Valid ipv4$ihl;
        meta.genv$optLen = tagged Valid genv$optLen;
        meta.ipv4$ttl = tagged Valid ipv4$ttl;
        meta.genv$oam = tagged Valid genv$oam;
        meta.genv$reserved2 = tagged Valid genv$reserved2;
        meta.genv$critical = tagged Valid genv$critical;
        meta.udp$srcPort = tagged Valid udp$srcPort;
        meta.genv$protoType = tagged Valid genv$protoType;
        meta.genv$ver = tagged Valid genv$ver;
        meta.udp$dstPort = tagged Valid udp$dstPort;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.ipv4$protocol = tagged Valid ipv4$protocol;
        meta.genv$reserved = tagged Valid genv$reserved;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv4GenvRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4NvgreRewriteRspT {pkt: .pkt, gre$s: .gre$s, ipv4$identification: .ipv4$identification, gre$R: .gre$R, nvgre$flow_id: .nvgre$flow_id, ipv4$ihl: .ipv4$ihl, gre$proto: .gre$proto, ipv4$ttl: .ipv4$ttl, gre$ver: .gre$ver, gre$S: .gre$S, gre$C: .gre$C, gre$recurse: .gre$recurse, nvgre$tni: .nvgre$tni, gre$K: .gre$K, gre$flags: .gre$flags, ethernet$etherType: .ethernet$etherType, ipv4$protocol: .ipv4$protocol, ipv4$version: .ipv4$version}: begin
        meta.gre$s = tagged Valid gre$s;
        meta.ipv4$identification = tagged Valid ipv4$identification;
        meta.gre$R = tagged Valid gre$R;
        meta.nvgre$flow_id = tagged Valid nvgre$flow_id;
        meta.ipv4$ihl = tagged Valid ipv4$ihl;
        meta.gre$proto = tagged Valid gre$proto;
        meta.ipv4$ttl = tagged Valid ipv4$ttl;
        meta.gre$ver = tagged Valid gre$ver;
        meta.gre$S = tagged Valid gre$S;
        meta.gre$C = tagged Valid gre$C;
        meta.gre$recurse = tagged Valid gre$recurse;
        meta.nvgre$tni = tagged Valid nvgre$tni;
        meta.gre$K = tagged Valid gre$K;
        meta.gre$flags = tagged Valid gre$flags;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.ipv4$protocol = tagged Valid ipv4$protocol;
        meta.ipv4$version = tagged Valid ipv4$version;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv4NvgreRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4GreRewriteRspT {pkt: .pkt, ipv4$protocol: .ipv4$protocol, ipv4$ihl: .ipv4$ihl, gre$proto: .gre$proto, ipv4$ttl: .ipv4$ttl, ipv4$identification: .ipv4$identification, ethernet$etherType: .ethernet$etherType, ipv4$version: .ipv4$version}: begin
        meta.ipv4$protocol = tagged Valid ipv4$protocol;
        meta.ipv4$ihl = tagged Valid ipv4$ihl;
        meta.gre$proto = tagged Valid gre$proto;
        meta.ipv4$ttl = tagged Valid ipv4$ttl;
        meta.ipv4$identification = tagged Valid ipv4$identification;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.ipv4$version = tagged Valid ipv4$version;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv4GreRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4IpRewriteRspT {pkt: .pkt, ipv4$protocol: .ipv4$protocol, ipv4$ihl: .ipv4$ihl, ipv4$ttl: .ipv4$ttl, ipv4$identification: .ipv4$identification, ethernet$etherType: .ethernet$etherType, ipv4$version: .ipv4$version}: begin
        meta.ipv4$protocol = tagged Valid ipv4$protocol;
        meta.ipv4$ihl = tagged Valid ipv4$ihl;
        meta.ipv4$ttl = tagged Valid ipv4$ttl;
        meta.ipv4$identification = tagged Valid ipv4$identification;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.ipv4$version = tagged Valid ipv4$version;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv4IpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv4ErspanT3RewriteRspT {pkt: .pkt, gre$S: .gre$S, ipv4$identification: .ipv4$identification, gre$s: .gre$s, ipv4$version: .ipv4$version, ipv4$ihl: .ipv4$ihl, gre$proto: .gre$proto, ipv4$ttl: .ipv4$ttl, gre$ver: .gre$ver, erspan_t3_header$timestamp: .erspan_t3_header$timestamp, gre$C: .gre$C, gre$recurse: .gre$recurse, erspan_t3_header$span_id: .erspan_t3_header$span_id, gre$K: .gre$K, erspan_t3_header$version: .erspan_t3_header$version, gre$flags: .gre$flags, erspan_t3_header$sgt_other: .erspan_t3_header$sgt_other, ipv4$protocol: .ipv4$protocol, gre$R: .gre$R}: begin
        meta.gre$S = tagged Valid gre$S;
        meta.ipv4$identification = tagged Valid ipv4$identification;
        meta.gre$s = tagged Valid gre$s;
        meta.ipv4$version = tagged Valid ipv4$version;
        meta.ipv4$ihl = tagged Valid ipv4$ihl;
        meta.gre$proto = tagged Valid gre$proto;
        meta.ipv4$ttl = tagged Valid ipv4$ttl;
        meta.gre$ver = tagged Valid gre$ver;
        meta.erspan_t3_header$timestamp = tagged Valid erspan_t3_header$timestamp;
        meta.gre$C = tagged Valid gre$C;
        meta.gre$recurse = tagged Valid gre$recurse;
        meta.erspan_t3_header$span_id = tagged Valid erspan_t3_header$span_id;
        meta.gre$K = tagged Valid gre$K;
        meta.erspan_t3_header$version = tagged Valid erspan_t3_header$version;
        meta.gre$flags = tagged Valid gre$flags;
        meta.erspan_t3_header$sgt_other = tagged Valid erspan_t3_header$sgt_other;
        meta.ipv4$protocol = tagged Valid ipv4$protocol;
        meta.gre$R = tagged Valid gre$R;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv4ErspanT3RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6GreRewriteRspT {pkt: .pkt, ipv6$version: .ipv6$version, ipv6$flowLabel: .ipv6$flowLabel, gre$proto: .gre$proto, ipv6$hopLimit: .ipv6$hopLimit, ipv6$trafficClass: .ipv6$trafficClass, ipv6$nextHdr: .ipv6$nextHdr, ethernet$etherType: .ethernet$etherType}: begin
        meta.ipv6$version = tagged Valid ipv6$version;
        meta.ipv6$flowLabel = tagged Valid ipv6$flowLabel;
        meta.gre$proto = tagged Valid gre$proto;
        meta.ipv6$hopLimit = tagged Valid ipv6$hopLimit;
        meta.ipv6$trafficClass = tagged Valid ipv6$trafficClass;
        meta.ipv6$nextHdr = tagged Valid ipv6$nextHdr;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv6GreRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6IpRewriteRspT {pkt: .pkt, ipv6$version: .ipv6$version, ipv6$payloadLen: .ipv6$payloadLen, ipv6$flowLabel: .ipv6$flowLabel, ipv6$hopLimit: .ipv6$hopLimit, ipv6$trafficClass: .ipv6$trafficClass, ipv6$nextHdr: .ipv6$nextHdr, ethernet$etherType: .ethernet$etherType}: begin
        meta.ipv6$version = tagged Valid ipv6$version;
        meta.ipv6$payloadLen = tagged Valid ipv6$payloadLen;
        meta.ipv6$flowLabel = tagged Valid ipv6$flowLabel;
        meta.ipv6$hopLimit = tagged Valid ipv6$hopLimit;
        meta.ipv6$trafficClass = tagged Valid ipv6$trafficClass;
        meta.ipv6$nextHdr = tagged Valid ipv6$nextHdr;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv6IpRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6NvgreRewriteRspT {pkt: .pkt, ipv6$version: .ipv6$version, gre$s: .gre$s, gre$R: .gre$R, nvgre$flow_id: .nvgre$flow_id, gre$proto: .gre$proto, gre$ver: .gre$ver, gre$S: .gre$S, ethernet$etherType: .ethernet$etherType, gre$C: .gre$C, gre$recurse: .gre$recurse, nvgre$tni: .nvgre$tni, ipv6$nextHdr: .ipv6$nextHdr, ipv6$flowLabel: .ipv6$flowLabel, gre$K: .gre$K, ipv6$trafficClass: .ipv6$trafficClass, gre$flags: .gre$flags, ipv6$hopLimit: .ipv6$hopLimit}: begin
        meta.ipv6$version = tagged Valid ipv6$version;
        meta.gre$s = tagged Valid gre$s;
        meta.gre$R = tagged Valid gre$R;
        meta.nvgre$flow_id = tagged Valid nvgre$flow_id;
        meta.gre$proto = tagged Valid gre$proto;
        meta.gre$ver = tagged Valid gre$ver;
        meta.gre$S = tagged Valid gre$S;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.gre$C = tagged Valid gre$C;
        meta.gre$recurse = tagged Valid gre$recurse;
        meta.nvgre$tni = tagged Valid nvgre$tni;
        meta.ipv6$nextHdr = tagged Valid ipv6$nextHdr;
        meta.ipv6$flowLabel = tagged Valid ipv6$flowLabel;
        meta.gre$K = tagged Valid gre$K;
        meta.ipv6$trafficClass = tagged Valid ipv6$trafficClass;
        meta.gre$flags = tagged Valid gre$flags;
        meta.ipv6$hopLimit = tagged Valid ipv6$hopLimit;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv6NvgreRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6VxlanRewriteRspT {pkt: .pkt, ipv6$version: .ipv6$version, udp$checksum: .udp$checksum, vxlan$vni: .vxlan$vni, vxlan$flags: .vxlan$flags, ipv6$nextHdr: .ipv6$nextHdr, vxlan$reserved2: .vxlan$reserved2, udp$srcPort: .udp$srcPort, ipv6$flowLabel: .ipv6$flowLabel, vxlan$reserved: .vxlan$reserved, ipv6$hopLimit: .ipv6$hopLimit, ipv6$trafficClass: .ipv6$trafficClass, udp$dstPort: .udp$dstPort, ethernet$etherType: .ethernet$etherType}: begin
        meta.ipv6$version = tagged Valid ipv6$version;
        meta.udp$checksum = tagged Valid udp$checksum;
        meta.vxlan$vni = tagged Valid vxlan$vni;
        meta.vxlan$flags = tagged Valid vxlan$flags;
        meta.ipv6$nextHdr = tagged Valid ipv6$nextHdr;
        meta.vxlan$reserved2 = tagged Valid vxlan$reserved2;
        meta.udp$srcPort = tagged Valid udp$srcPort;
        meta.ipv6$flowLabel = tagged Valid ipv6$flowLabel;
        meta.vxlan$reserved = tagged Valid vxlan$reserved;
        meta.ipv6$hopLimit = tagged Valid ipv6$hopLimit;
        meta.ipv6$trafficClass = tagged Valid ipv6$trafficClass;
        meta.udp$dstPort = tagged Valid udp$dstPort;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv6VxlanRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6GenvRewriteRspT {pkt: .pkt, genv$vni: .genv$vni, ipv6$trafficClass: .ipv6$trafficClass, udp$checksum: .udp$checksum, ipv6$version: .ipv6$version, genv$optLen: .genv$optLen, ipv6$nextHdr: .ipv6$nextHdr, genv$oam: .genv$oam, genv$reserved2: .genv$reserved2, ethernet$etherType: .ethernet$etherType, genv$critical: .genv$critical, udp$srcPort: .udp$srcPort, ipv6$flowLabel: .ipv6$flowLabel, genv$protoType: .genv$protoType, genv$ver: .genv$ver, udp$dstPort: .udp$dstPort, ipv6$hopLimit: .ipv6$hopLimit, genv$reserved: .genv$reserved}: begin
        meta.genv$vni = tagged Valid genv$vni;
        meta.ipv6$trafficClass = tagged Valid ipv6$trafficClass;
        meta.udp$checksum = tagged Valid udp$checksum;
        meta.ipv6$version = tagged Valid ipv6$version;
        meta.genv$optLen = tagged Valid genv$optLen;
        meta.ipv6$nextHdr = tagged Valid ipv6$nextHdr;
        meta.genv$oam = tagged Valid genv$oam;
        meta.genv$reserved2 = tagged Valid genv$reserved2;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.genv$critical = tagged Valid genv$critical;
        meta.udp$srcPort = tagged Valid udp$srcPort;
        meta.ipv6$flowLabel = tagged Valid ipv6$flowLabel;
        meta.genv$protoType = tagged Valid genv$protoType;
        meta.genv$ver = tagged Valid genv$ver;
        meta.udp$dstPort = tagged Valid udp$dstPort;
        meta.ipv6$hopLimit = tagged Valid ipv6$hopLimit;
        meta.genv$reserved = tagged Valid genv$reserved;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv6GenvRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged Ipv6ErspanT3RewriteRspT {pkt: .pkt, ipv6$version: .ipv6$version, gre$S: .gre$S, ipv6$trafficClass: .ipv6$trafficClass, gre$s: .gre$s, ipv6$hopLimit: .ipv6$hopLimit, ipv6$flowLabel: .ipv6$flowLabel, gre$proto: .gre$proto, gre$ver: .gre$ver, erspan_t3_header$timestamp: .erspan_t3_header$timestamp, gre$C: .gre$C, gre$recurse: .gre$recurse, ipv6$nextHdr: .ipv6$nextHdr, erspan_t3_header$span_id: .erspan_t3_header$span_id, gre$K: .gre$K, erspan_t3_header$version: .erspan_t3_header$version, gre$flags: .gre$flags, erspan_t3_header$sgt_other: .erspan_t3_header$sgt_other, gre$R: .gre$R}: begin
        meta.ipv6$version = tagged Valid ipv6$version;
        meta.gre$S = tagged Valid gre$S;
        meta.ipv6$trafficClass = tagged Valid ipv6$trafficClass;
        meta.gre$s = tagged Valid gre$s;
        meta.ipv6$hopLimit = tagged Valid ipv6$hopLimit;
        meta.ipv6$flowLabel = tagged Valid ipv6$flowLabel;
        meta.gre$proto = tagged Valid gre$proto;
        meta.gre$ver = tagged Valid gre$ver;
        meta.erspan_t3_header$timestamp = tagged Valid erspan_t3_header$timestamp;
        meta.gre$C = tagged Valid gre$C;
        meta.gre$recurse = tagged Valid gre$recurse;
        meta.ipv6$nextHdr = tagged Valid ipv6$nextHdr;
        meta.erspan_t3_header$span_id = tagged Valid erspan_t3_header$span_id;
        meta.gre$K = tagged Valid gre$K;
        meta.erspan_t3_header$version = tagged Valid erspan_t3_header$version;
        meta.gre$flags = tagged Valid gre$flags;
        meta.erspan_t3_header$sgt_other = tagged Valid erspan_t3_header$sgt_other;
        meta.gre$R = tagged Valid gre$R;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterIpv6ErspanT3RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MplsEthernetPush1RewriteRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterMplsEthernetPush1RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MplsIpPush1RewriteRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterMplsIpPush1RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MplsEthernetPush2RewriteRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterMplsEthernetPush2RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MplsIpPush2RewriteRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterMplsIpPush2RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MplsEthernetPush3RewriteRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterMplsEthernetPush3RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged MplsIpPush3RewriteRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterMplsIpPush3RewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FabricRewriteRspT {pkt: .pkt, tunnel_metadata$tunnel_index: .tunnel_metadata$tunnel_index}: begin
        meta.tunnel_metadata$tunnel_index = tagged Valid tunnel_metadata$tunnel_index;
        MetadataResponse rsp = tagged TunnelEncapProcessOuterFabricRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
  interface next_control_state_8 = toClient(bbReqFifo[8], bbRspFifo[8]);
  interface next_control_state_9 = toClient(bbReqFifo[9], bbRspFifo[9]);
  interface next_control_state_10 = toClient(bbReqFifo[10], bbRspFifo[10]);
  interface next_control_state_11 = toClient(bbReqFifo[11], bbRspFifo[11]);
  interface next_control_state_12 = toClient(bbReqFifo[12], bbRspFifo[12]);
  interface next_control_state_13 = toClient(bbReqFifo[13], bbRspFifo[13]);
  interface next_control_state_14 = toClient(bbReqFifo[14], bbRspFifo[14]);
  interface next_control_state_15 = toClient(bbReqFifo[15], bbRspFifo[15]);
  interface next_control_state_16 = toClient(bbReqFifo[16], bbRspFifo[16]);
  interface next_control_state_17 = toClient(bbReqFifo[17], bbRspFifo[17]);
  interface next_control_state_18 = toClient(bbReqFifo[18], bbRspFifo[18]);
  interface next_control_state_19 = toClient(bbReqFifo[19], bbRspFifo[19]);
endmodule

// ====== TUNNEL_MTU ======

typedef struct {
  Bit#(4) padding;
  Bit#(14) tunnel_metadata$tunnel_index;
} TunnelMtuReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_MTU,
  TUNNEL_MTU_CHECK,
  TUNNEL_MTU_MISS
} TunnelMtuActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelMtuActionT _action;
  Bit#(16) runtime_l3_mtu;
} TunnelMtuRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(18)) matchtable_read_tunnel_mtu(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_tunnel_mtu(Bit#(18) msgtype, Bit#(18) data);
`endif
instance MatchTableSim#(92, 18, 18);
  function ActionValue#(Bit#(18)) matchtable_read(Bit#(92) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_tunnel_mtu(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(92) id, Bit#(18) key, Bit#(18) data);
    action
      matchtable_write_tunnel_mtu(key, data);
    endaction
  endfunction

endinstance
interface TunnelMtu;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkTunnelMtu  (TunnelMtu);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(92, 1024, SizeOf#(TunnelMtuReqT), SizeOf#(TunnelMtuRspT)) matchTable <- mkMatchTable("tunnel_mtu.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$tunnel_index = fromMaybe(?, meta.tunnel_metadata$tunnel_index);
    TunnelMtuReqT req = TunnelMtuReqT {tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelMtuRspT resp = unpack(data);
      case (resp._action) matches
        TUNNEL_MTU_CHECK: begin
          BBRequest req = tagged TunnelMtuCheckReqT {pkt: pkt, runtime_l3_mtu: resp.runtime_l3_mtu};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        TUNNEL_MTU_MISS: begin
          BBRequest req = tagged TunnelMtuMissReqT {pkt: pkt};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged TunnelMtuCheckRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelMtuTunnelMtuCheckRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged TunnelMtuMissRspT {pkt: .pkt, l3_metadata$l3_mtu_check: .l3_metadata$l3_mtu_check}: begin
        meta.l3_metadata$l3_mtu_check = tagged Valid l3_metadata$l3_mtu_check;
        MetadataResponse rsp = tagged TunnelMtuTunnelMtuMissRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== TUNNEL_REWRITE ======

typedef struct {
  Bit#(4) padding;
  Bit#(14) tunnel_metadata$tunnel_index;
} TunnelRewriteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_REWRITE,
  NOP,
  SET_TUNNEL_REWRITE_DETAILS,
  SET_MPLS_REWRITE_PUSH1,
  SET_MPLS_REWRITE_PUSH2,
  SET_MPLS_REWRITE_PUSH3,
  CPU_RX_REWRITE,
  FABRIC_UNICAST_REWRITE,
  FABRIC_MULTICAST_REWRITE
} TunnelRewriteActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelRewriteActionT _action;
  Bit#(16) runtime_outer_bd;
  Bit#(9) runtime_smac_idx;
  Bit#(14) runtime_dmac_idx;
  Bit#(9) runtime_sip_index;
  Bit#(14) runtime_dip_index;
  Bit#(20) runtime_label1;
  Bit#(3) runtime_exp1;
  Bit#(8) runtime_ttl1;
  Bit#(20) runtime_label2;
  Bit#(3) runtime_exp2;
  Bit#(8) runtime_ttl2;
  Bit#(20) runtime_label3;
  Bit#(3) runtime_exp3;
  Bit#(8) runtime_ttl3;
  Bit#(16) runtime_fabric_mgid;
} TunnelRewriteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(175)) matchtable_read_tunnel_rewrite(Bit#(18) msgtype);
import "BDPI" function Action matchtable_write_tunnel_rewrite(Bit#(18) msgtype, Bit#(175) data);
`endif
instance MatchTableSim#(91, 18, 175);
  function ActionValue#(Bit#(175)) matchtable_read(Bit#(91) id, Bit#(18) key);
    actionvalue
      let v <- matchtable_read_tunnel_rewrite(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(91) id, Bit#(18) key, Bit#(175) data);
    action
      matchtable_write_tunnel_rewrite(key, data);
    endaction
  endfunction

endinstance
interface TunnelRewrite;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
  interface Client #(BBRequest, BBResponse) next_control_state_3;
  interface Client #(BBRequest, BBResponse) next_control_state_4;
  interface Client #(BBRequest, BBResponse) next_control_state_5;
  interface Client #(BBRequest, BBResponse) next_control_state_6;
  interface Client #(BBRequest, BBResponse) next_control_state_7;
endinterface
(* synthesize *)
module mkTunnelRewrite  (TunnelRewrite);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(8, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(8, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(91, 1024, SizeOf#(TunnelRewriteReqT), SizeOf#(TunnelRewriteRspT)) matchTable <- mkMatchTable("tunnel_rewrite.dat");
  Vector#(8, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(8) readyChannel = -1;
  for (Integer i=7; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$tunnel_index = fromMaybe(?, meta.tunnel_metadata$tunnel_index);
    TunnelRewriteReqT req = TunnelRewriteReqT {tunnel_metadata$tunnel_index: tunnel_metadata$tunnel_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelRewriteRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        SET_TUNNEL_REWRITE_DETAILS: begin
          BBRequest req = tagged SetTunnelRewriteDetailsReqT {pkt: pkt, runtime_outer_bd: resp.runtime_outer_bd, runtime_sip_index: resp.runtime_sip_index, runtime_dip_index: resp.runtime_dip_index, runtime_dmac_idx: resp.runtime_dmac_idx, runtime_smac_idx: resp.runtime_smac_idx};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        SET_MPLS_REWRITE_PUSH1: begin
          BBRequest req = tagged SetMplsRewritePush1ReqT {pkt: pkt, runtime_ttl1: resp.runtime_ttl1, runtime_exp1: resp.runtime_exp1, runtime_label1: resp.runtime_label1, runtime_dmac_idx: resp.runtime_dmac_idx, runtime_smac_idx: resp.runtime_smac_idx};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
        SET_MPLS_REWRITE_PUSH2: begin
          BBRequest req = tagged SetMplsRewritePush2ReqT {pkt: pkt, runtime_exp1: resp.runtime_exp1, runtime_ttl2: resp.runtime_ttl2, runtime_smac_idx: resp.runtime_smac_idx, runtime_ttl1: resp.runtime_ttl1, runtime_label2: resp.runtime_label2, runtime_exp2: resp.runtime_exp2, runtime_label1: resp.runtime_label1, runtime_dmac_idx: resp.runtime_dmac_idx};
          bbReqFifo[3].enq(req); //FIXME: replace with RXTX.
        end
        SET_MPLS_REWRITE_PUSH3: begin
          BBRequest req = tagged SetMplsRewritePush3ReqT {pkt: pkt, runtime_exp3: resp.runtime_exp3, runtime_exp1: resp.runtime_exp1, runtime_ttl2: resp.runtime_ttl2, runtime_label3: resp.runtime_label3, runtime_ttl1: resp.runtime_ttl1, runtime_label2: resp.runtime_label2, runtime_exp2: resp.runtime_exp2, runtime_label1: resp.runtime_label1, runtime_smac_idx: resp.runtime_smac_idx, runtime_ttl3: resp.runtime_ttl3, runtime_dmac_idx: resp.runtime_dmac_idx};
          bbReqFifo[4].enq(req); //FIXME: replace with RXTX.
        end
        CPU_RX_REWRITE: begin
          BBRequest req = tagged CpuRxRewriteReqT {pkt: pkt, ingress_metadata$bd: ingress_metadata$bd, fabric_metadata$reason_code: fabric_metadata$reason_code, ingress_metadata$ingress_port: ingress_metadata$ingress_port, ingress_metadata$ifindex: ingress_metadata$ifindex, ethernet$etherType: ethernet$etherType};
          bbReqFifo[5].enq(req); //FIXME: replace with RXTX.
        end
        FABRIC_UNICAST_REWRITE: begin
          BBRequest req = tagged FabricUnicastRewriteReqT {pkt: pkt, l3_metadata$nexthop_index: l3_metadata$nexthop_index, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type, l3_metadata$routed: l3_metadata$routed, fabric_metadata$dst_device: fabric_metadata$dst_device, fabric_metadata$dst_port: fabric_metadata$dst_port, ethernet$etherType: ethernet$etherType, l3_metadata$outer_routed: l3_metadata$outer_routed};
          bbReqFifo[6].enq(req); //FIXME: replace with RXTX.
        end
        FABRIC_MULTICAST_REWRITE: begin
          BBRequest req = tagged FabricMulticastRewriteReqT {pkt: pkt, multicast_metadata$mcast_grp: multicast_metadata$mcast_grp, ingress_metadata$bd: ingress_metadata$bd, tunnel_metadata$ingress_tunnel_type: tunnel_metadata$ingress_tunnel_type, l3_metadata$routed: l3_metadata$routed, tunnel_metadata$tunnel_terminate: tunnel_metadata$tunnel_terminate, ingress_metadata$ifindex: ingress_metadata$ifindex, ethernet$etherType: ethernet$etherType, l3_metadata$outer_routed: l3_metadata$outer_routed, runtime_fabric_mgid: resp.runtime_fabric_mgid};
          bbReqFifo[7].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelRewriteNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetTunnelRewriteDetailsRspT {pkt: .pkt, egress_metadata$outer_bd: .egress_metadata$outer_bd, tunnel_metadata$tunnel_src_index: .tunnel_metadata$tunnel_src_index, tunnel_metadata$tunnel_dst_index: .tunnel_metadata$tunnel_dst_index, tunnel_metadata$tunnel_dmac_index: .tunnel_metadata$tunnel_dmac_index, tunnel_metadata$tunnel_smac_index: .tunnel_metadata$tunnel_smac_index}: begin
        meta.egress_metadata$outer_bd = tagged Valid egress_metadata$outer_bd;
        meta.tunnel_metadata$tunnel_src_index = tagged Valid tunnel_metadata$tunnel_src_index;
        meta.tunnel_metadata$tunnel_dst_index = tagged Valid tunnel_metadata$tunnel_dst_index;
        meta.tunnel_metadata$tunnel_dmac_index = tagged Valid tunnel_metadata$tunnel_dmac_index;
        meta.tunnel_metadata$tunnel_smac_index = tagged Valid tunnel_metadata$tunnel_smac_index;
        MetadataResponse rsp = tagged TunnelRewriteSetTunnelRewriteDetailsRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMplsRewritePush1RspT {pkt: .pkt, tunnel_metadata$tunnel_smac_index: .tunnel_metadata$tunnel_smac_index, mpls0$exp: .mpls0$exp, mpls0$ttl: .mpls0$ttl, mpls0$bos: .mpls0$bos, tunnel_metadata$tunnel_dmac_index: .tunnel_metadata$tunnel_dmac_index, mpls0$label: .mpls0$label}: begin
        meta.tunnel_metadata$tunnel_smac_index = tagged Valid tunnel_metadata$tunnel_smac_index;
        meta.mpls0$exp = tagged Valid mpls0$exp;
        meta.mpls0$ttl = tagged Valid mpls0$ttl;
        meta.mpls0$bos = tagged Valid mpls0$bos;
        meta.tunnel_metadata$tunnel_dmac_index = tagged Valid tunnel_metadata$tunnel_dmac_index;
        meta.mpls0$label = tagged Valid mpls0$label;
        MetadataResponse rsp = tagged TunnelRewriteSetMplsRewritePush1RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMplsRewritePush2RspT {pkt: .pkt, mpls1$ttl: .mpls1$ttl, tunnel_metadata$tunnel_smac_index: .tunnel_metadata$tunnel_smac_index, mpls1$exp: .mpls1$exp, mpls0$exp: .mpls0$exp, mpls0$ttl: .mpls0$ttl, mpls1$label: .mpls1$label, mpls0$bos: .mpls0$bos, mpls1$bos: .mpls1$bos, tunnel_metadata$tunnel_dmac_index: .tunnel_metadata$tunnel_dmac_index, mpls0$label: .mpls0$label}: begin
        meta.mpls1$ttl = tagged Valid mpls1$ttl;
        meta.tunnel_metadata$tunnel_smac_index = tagged Valid tunnel_metadata$tunnel_smac_index;
        meta.mpls1$exp = tagged Valid mpls1$exp;
        meta.mpls0$exp = tagged Valid mpls0$exp;
        meta.mpls0$ttl = tagged Valid mpls0$ttl;
        meta.mpls1$label = tagged Valid mpls1$label;
        meta.mpls0$bos = tagged Valid mpls0$bos;
        meta.mpls1$bos = tagged Valid mpls1$bos;
        meta.tunnel_metadata$tunnel_dmac_index = tagged Valid tunnel_metadata$tunnel_dmac_index;
        meta.mpls0$label = tagged Valid mpls0$label;
        MetadataResponse rsp = tagged TunnelRewriteSetMplsRewritePush2RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged SetMplsRewritePush3RspT {pkt: .pkt, mpls1$ttl: .mpls1$ttl, mpls1$exp: .mpls1$exp, mpls2$bos: .mpls2$bos, tunnel_metadata$tunnel_smac_index: .tunnel_metadata$tunnel_smac_index, mpls1$label: .mpls1$label, mpls0$bos: .mpls0$bos, mpls2$exp: .mpls2$exp, mpls2$ttl: .mpls2$ttl, mpls0$exp: .mpls0$exp, tunnel_metadata$tunnel_dmac_index: .tunnel_metadata$tunnel_dmac_index, mpls0$ttl: .mpls0$ttl, mpls2$label: .mpls2$label, mpls1$bos: .mpls1$bos, mpls0$label: .mpls0$label}: begin
        meta.mpls1$ttl = tagged Valid mpls1$ttl;
        meta.mpls1$exp = tagged Valid mpls1$exp;
        meta.mpls2$bos = tagged Valid mpls2$bos;
        meta.tunnel_metadata$tunnel_smac_index = tagged Valid tunnel_metadata$tunnel_smac_index;
        meta.mpls1$label = tagged Valid mpls1$label;
        meta.mpls0$bos = tagged Valid mpls0$bos;
        meta.mpls2$exp = tagged Valid mpls2$exp;
        meta.mpls2$ttl = tagged Valid mpls2$ttl;
        meta.mpls0$exp = tagged Valid mpls0$exp;
        meta.tunnel_metadata$tunnel_dmac_index = tagged Valid tunnel_metadata$tunnel_dmac_index;
        meta.mpls0$ttl = tagged Valid mpls0$ttl;
        meta.mpls2$label = tagged Valid mpls2$label;
        meta.mpls1$bos = tagged Valid mpls1$bos;
        meta.mpls0$label = tagged Valid mpls0$label;
        MetadataResponse rsp = tagged TunnelRewriteSetMplsRewritePush3RspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged CpuRxRewriteRspT {pkt: .pkt, fabric_header$packetType: .fabric_header$packetType, fabric_header_cpu$reasonCode: .fabric_header_cpu$reasonCode, fabric_header_cpu$ingressPort: .fabric_header_cpu$ingressPort, fabric_header_cpu$ingressIfindex: .fabric_header_cpu$ingressIfindex, fabric_payload_header$etherType: .fabric_payload_header$etherType, fabric_header_cpu$ingressBd: .fabric_header_cpu$ingressBd, fabric_header$headerVersion: .fabric_header$headerVersion, fabric_header$packetVersion: .fabric_header$packetVersion, ethernet$etherType: .ethernet$etherType, fabric_header$pad1: .fabric_header$pad1}: begin
        meta.fabric_header$packetType = tagged Valid fabric_header$packetType;
        meta.fabric_header_cpu$reasonCode = tagged Valid fabric_header_cpu$reasonCode;
        meta.fabric_header_cpu$ingressPort = tagged Valid fabric_header_cpu$ingressPort;
        meta.fabric_header_cpu$ingressIfindex = tagged Valid fabric_header_cpu$ingressIfindex;
        meta.fabric_payload_header$etherType = tagged Valid fabric_payload_header$etherType;
        meta.fabric_header_cpu$ingressBd = tagged Valid fabric_header_cpu$ingressBd;
        meta.fabric_header$headerVersion = tagged Valid fabric_header$headerVersion;
        meta.fabric_header$packetVersion = tagged Valid fabric_header$packetVersion;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.fabric_header$pad1 = tagged Valid fabric_header$pad1;
        MetadataResponse rsp = tagged TunnelRewriteCpuRxRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FabricUnicastRewriteRspT {pkt: .pkt, fabric_header$packetType: .fabric_header$packetType, fabric_header_unicast$outerRouted: .fabric_header_unicast$outerRouted, fabric_header_unicast$tunnelTerminate: .fabric_header_unicast$tunnelTerminate, fabric_payload_header$etherType: .fabric_payload_header$etherType, fabric_header$dstDevice: .fabric_header$dstDevice, fabric_header_unicast$ingressTunnelType: .fabric_header_unicast$ingressTunnelType, fabric_header$dstPortOrGroup: .fabric_header$dstPortOrGroup, fabric_header_unicast$nexthopIndex: .fabric_header_unicast$nexthopIndex, fabric_header_unicast$routed: .fabric_header_unicast$routed, fabric_header$pad1: .fabric_header$pad1, fabric_header$packetVersion: .fabric_header$packetVersion, ethernet$etherType: .ethernet$etherType, fabric_header$headerVersion: .fabric_header$headerVersion}: begin
        meta.fabric_header$packetType = tagged Valid fabric_header$packetType;
        meta.fabric_header_unicast$outerRouted = tagged Valid fabric_header_unicast$outerRouted;
        meta.fabric_header_unicast$tunnelTerminate = tagged Valid fabric_header_unicast$tunnelTerminate;
        meta.fabric_payload_header$etherType = tagged Valid fabric_payload_header$etherType;
        meta.fabric_header$dstDevice = tagged Valid fabric_header$dstDevice;
        meta.fabric_header_unicast$ingressTunnelType = tagged Valid fabric_header_unicast$ingressTunnelType;
        meta.fabric_header$dstPortOrGroup = tagged Valid fabric_header$dstPortOrGroup;
        meta.fabric_header_unicast$nexthopIndex = tagged Valid fabric_header_unicast$nexthopIndex;
        meta.fabric_header_unicast$routed = tagged Valid fabric_header_unicast$routed;
        meta.fabric_header$pad1 = tagged Valid fabric_header$pad1;
        meta.fabric_header$packetVersion = tagged Valid fabric_header$packetVersion;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.fabric_header$headerVersion = tagged Valid fabric_header$headerVersion;
        MetadataResponse rsp = tagged TunnelRewriteFabricUnicastRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged FabricMulticastRewriteRspT {pkt: .pkt, fabric_header$packetType: .fabric_header$packetType, fabric_header_multicast$tunnelTerminate: .fabric_header_multicast$tunnelTerminate, fabric_header_multicast$routed: .fabric_header_multicast$routed, fabric_header_multicast$ingressTunnelType: .fabric_header_multicast$ingressTunnelType, fabric_header$dstDevice: .fabric_header$dstDevice, fabric_header_multicast$outerRouted: .fabric_header_multicast$outerRouted, fabric_header_multicast$ingressIfindex: .fabric_header_multicast$ingressIfindex, fabric_header$dstPortOrGroup: .fabric_header$dstPortOrGroup, fabric_payload_header$etherType: .fabric_payload_header$etherType, fabric_header_multicast$ingressBd: .fabric_header_multicast$ingressBd, fabric_header_multicast$mcastGrp: .fabric_header_multicast$mcastGrp, fabric_header$pad1: .fabric_header$pad1, fabric_header$packetVersion: .fabric_header$packetVersion, ethernet$etherType: .ethernet$etherType, fabric_header$headerVersion: .fabric_header$headerVersion}: begin
        meta.fabric_header$packetType = tagged Valid fabric_header$packetType;
        meta.fabric_header_multicast$tunnelTerminate = tagged Valid fabric_header_multicast$tunnelTerminate;
        meta.fabric_header_multicast$routed = tagged Valid fabric_header_multicast$routed;
        meta.fabric_header_multicast$ingressTunnelType = tagged Valid fabric_header_multicast$ingressTunnelType;
        meta.fabric_header$dstDevice = tagged Valid fabric_header$dstDevice;
        meta.fabric_header_multicast$outerRouted = tagged Valid fabric_header_multicast$outerRouted;
        meta.fabric_header_multicast$ingressIfindex = tagged Valid fabric_header_multicast$ingressIfindex;
        meta.fabric_header$dstPortOrGroup = tagged Valid fabric_header$dstPortOrGroup;
        meta.fabric_payload_header$etherType = tagged Valid fabric_payload_header$etherType;
        meta.fabric_header_multicast$ingressBd = tagged Valid fabric_header_multicast$ingressBd;
        meta.fabric_header_multicast$mcastGrp = tagged Valid fabric_header_multicast$mcastGrp;
        meta.fabric_header$pad1 = tagged Valid fabric_header$pad1;
        meta.fabric_header$packetVersion = tagged Valid fabric_header$packetVersion;
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        meta.fabric_header$headerVersion = tagged Valid fabric_header$headerVersion;
        MetadataResponse rsp = tagged TunnelRewriteFabricMulticastRewriteRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
  interface next_control_state_3 = toClient(bbReqFifo[3], bbRspFifo[3]);
  interface next_control_state_4 = toClient(bbReqFifo[4], bbRspFifo[4]);
  interface next_control_state_5 = toClient(bbReqFifo[5], bbRspFifo[5]);
  interface next_control_state_6 = toClient(bbReqFifo[6], bbRspFifo[6]);
  interface next_control_state_7 = toClient(bbReqFifo[7], bbRspFifo[7]);
endmodule

// ====== TUNNEL_SMAC_REWRITE ======

typedef struct {
  Bit#(9) tunnel_metadata$tunnel_smac_index;
} TunnelSmacRewriteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_SMAC_REWRITE,
  NOP,
  REWRITE_TUNNEL_SMAC
} TunnelSmacRewriteActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelSmacRewriteActionT _action;
  Bit#(48) runtime_smac;
} TunnelSmacRewriteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(50)) matchtable_read_tunnel_smac_rewrite(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_tunnel_smac_rewrite(Bit#(9) msgtype, Bit#(50) data);
`endif
instance MatchTableSim#(95, 9, 50);
  function ActionValue#(Bit#(50)) matchtable_read(Bit#(95) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_tunnel_smac_rewrite(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(95) id, Bit#(9) key, Bit#(50) data);
    action
      matchtable_write_tunnel_smac_rewrite(key, data);
    endaction
  endfunction

endinstance
interface TunnelSmacRewrite;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
endinterface
(* synthesize *)
module mkTunnelSmacRewrite  (TunnelSmacRewrite);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(2, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(2, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(95, 1024, SizeOf#(TunnelSmacRewriteReqT), SizeOf#(TunnelSmacRewriteRspT)) matchTable <- mkMatchTable("tunnel_smac_rewrite.dat");
  Vector#(2, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(2) readyChannel = -1;
  for (Integer i=1; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$tunnel_smac_index = fromMaybe(?, meta.tunnel_metadata$tunnel_smac_index);
    TunnelSmacRewriteReqT req = TunnelSmacRewriteReqT {tunnel_metadata$tunnel_smac_index: tunnel_metadata$tunnel_smac_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelSmacRewriteRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        REWRITE_TUNNEL_SMAC: begin
          BBRequest req = tagged RewriteTunnelSmacReqT {pkt: pkt, runtime_smac: resp.runtime_smac};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelSmacRewriteNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RewriteTunnelSmacRspT {pkt: .pkt, ethernet$srcAddr: .ethernet$srcAddr}: begin
        meta.ethernet$srcAddr = tagged Valid ethernet$srcAddr;
        MetadataResponse rsp = tagged TunnelSmacRewriteRewriteTunnelSmacRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
endmodule

// ====== TUNNEL_SRC_REWRITE ======

typedef struct {
  Bit#(9) tunnel_metadata$tunnel_src_index;
} TunnelSrcRewriteReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_TUNNEL_SRC_REWRITE,
  NOP,
  REWRITE_TUNNEL_IPV4_SRC,
  REWRITE_TUNNEL_IPV6_SRC
} TunnelSrcRewriteActionT deriving (Bits, Eq, FShow);
typedef struct {
  TunnelSrcRewriteActionT _action;
  Bit#(32) runtime_ip;
} TunnelSrcRewriteRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(34)) matchtable_read_tunnel_src_rewrite(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_tunnel_src_rewrite(Bit#(9) msgtype, Bit#(34) data);
`endif
instance MatchTableSim#(93, 9, 34);
  function ActionValue#(Bit#(34)) matchtable_read(Bit#(93) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_tunnel_src_rewrite(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(93) id, Bit#(9) key, Bit#(34) data);
    action
      matchtable_write_tunnel_src_rewrite(key, data);
    endaction
  endfunction

endinstance
interface TunnelSrcRewrite;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkTunnelSrcRewrite  (TunnelSrcRewrite);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(93, 1024, SizeOf#(TunnelSrcRewriteReqT), SizeOf#(TunnelSrcRewriteRspT)) matchTable <- mkMatchTable("tunnel_src_rewrite.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let tunnel_metadata$tunnel_src_index = fromMaybe(?, meta.tunnel_metadata$tunnel_src_index);
    TunnelSrcRewriteReqT req = TunnelSrcRewriteReqT {tunnel_metadata$tunnel_src_index: tunnel_metadata$tunnel_src_index};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      TunnelSrcRewriteRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        REWRITE_TUNNEL_IPV4_SRC: begin
          BBRequest req = tagged RewriteTunnelIpv4SrcReqT {pkt: pkt, runtime_ip: resp.runtime_ip};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        REWRITE_TUNNEL_IPV6_SRC: begin
          BBRequest req = tagged RewriteTunnelIpv6SrcReqT {pkt: pkt, runtime_ip: resp.runtime_ip};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged TunnelSrcRewriteNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RewriteTunnelIpv4SrcRspT {pkt: .pkt, ipv4$srcAddr: .ipv4$srcAddr}: begin
        meta.ipv4$srcAddr = tagged Valid ipv4$srcAddr;
        MetadataResponse rsp = tagged TunnelSrcRewriteRewriteTunnelIpv4SrcRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RewriteTunnelIpv6SrcRspT {pkt: .pkt, ipv6$srcAddr: .ipv6$srcAddr}: begin
        meta.ipv6$srcAddr = tagged Valid ipv6$srcAddr;
        MetadataResponse rsp = tagged TunnelSrcRewriteRewriteTunnelIpv6SrcRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== VLAN_DECAP ======

typedef struct {
  Bit#(7) padding;
  Bit#(Bool) valid_vlan_tag_0;
  Bit#(Bool) valid_vlan_tag_1;
} VlanDecapReqT deriving (Bits, Eq, FShow);
typedef enum {
  DEFAULT_VLAN_DECAP,
  NOP,
  REMOVE_VLAN_SINGLE_TAGGED,
  REMOVE_VLAN_DOUBLE_TAGGED
} VlanDecapActionT deriving (Bits, Eq, FShow);
typedef struct {
  VlanDecapActionT _action;
} VlanDecapRspT deriving (Bits, Eq, FShow);
`ifndef SVDPI
import "BDPI" function ActionValue#(Bit#(2)) matchtable_read_vlan_decap(Bit#(9) msgtype);
import "BDPI" function Action matchtable_write_vlan_decap(Bit#(9) msgtype, Bit#(2) data);
`endif
instance MatchTableSim#(82, 9, 2);
  function ActionValue#(Bit#(2)) matchtable_read(Bit#(82) id, Bit#(9) key);
    actionvalue
      let v <- matchtable_read_vlan_decap(key);
      return v;
    endactionvalue
  endfunction

  function Action matchtable_write(Bit#(82) id, Bit#(9) key, Bit#(2) data);
    action
      matchtable_write_vlan_decap(key, data);
    endaction
  endfunction

endinstance
interface VlanDecap;
  interface Server #(MetadataRequest, MetadataResponse) prev_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_0;
  interface Client #(BBRequest, BBResponse) next_control_state_1;
  interface Client #(BBRequest, BBResponse) next_control_state_2;
endinterface
(* synthesize *)
module mkVlanDecap  (VlanDecap);
  RX #(MetadataRequest) rx_metadata <- mkRX;
  let rx_info_metadata = rx_metadata.u;
  TX #(MetadataResponse) tx_metadata <- mkTX;
  let tx_info_metadata = tx_metadata.u;
  Vector#(3, FIFOF#(BBRequest)) bbReqFifo <- replicateM(mkFIFOF);
  Vector#(3, FIFOF#(BBResponse)) bbRspFifo <- replicateM(mkFIFOF);
  FIFOF#(PacketInstance) packet_ff <- mkFIFOF;
  MatchTable#(82, 1024, SizeOf#(VlanDecapReqT), SizeOf#(VlanDecapRspT)) matchTable <- mkMatchTable("vlan_decap.dat");
  Vector#(3, Bool) readyBits = map(fifoNotEmpty, bbRspFifo);
  Bool interruptStatus = False;
  Bit#(3) readyChannel = -1;
  for (Integer i=2; i>=0; i=i-1) begin
      if (readyBits[i]) begin
          interruptStatus = True;
          readyChannel = fromInteger(i);
      end
  end

  Vector#(2, FIFOF#(MetadataT)) metadata_ff <- replicateM(mkFIFOF);
  rule rl_handle_request;
    let data = rx_info_metadata.first;
    rx_info_metadata.deq;
    let meta = data.meta;
    let pkt = data.pkt;
    let v$l$a$n$_$t$a$g$_$$0$ = fromMaybe(?, meta.v$l$a$n$_$t$a$g$_$$0$);
    let v$l$a$n$_$t$a$g$_$$1$ = fromMaybe(?, meta.v$l$a$n$_$t$a$g$_$$1$);
    VlanDecapReqT req = VlanDecapReqT {v$l$a$n$_$t$a$g$_$$0$: v$l$a$n$_$t$a$g$_$$0$,v$l$a$n$_$t$a$g$_$$1$: v$l$a$n$_$t$a$g$_$$1$};
    matchTable.lookupPort.request.put(pack(req));
    packet_ff.enq(pkt);
    metadata_ff[0].enq(meta);
  endrule

  rule rl_handle_execute;
    let rsp <- matchTable.lookupPort.response.get;
    let pkt <- toGet(packet_ff).get;
    let meta <- toGet(metadata_ff[0]).get;
    if (rsp matches tagged Valid .data) begin
      VlanDecapRspT resp = unpack(data);
      case (resp._action) matches
        NOP: begin
          BBRequest req = tagged NopReqT {pkt: pkt};
          bbReqFifo[0].enq(req); //FIXME: replace with RXTX.
        end
        REMOVE_VLAN_SINGLE_TAGGED: begin
          BBRequest req = tagged RemoveVlanSingleTaggedReqT {pkt: pkt, vlan_tag_0$etherType: vlan_tag_0$etherType};
          bbReqFifo[1].enq(req); //FIXME: replace with RXTX.
        end
        REMOVE_VLAN_DOUBLE_TAGGED: begin
          BBRequest req = tagged RemoveVlanDoubleTaggedReqT {pkt: pkt, vlan_tag_1$etherType: vlan_tag_1$etherType};
          bbReqFifo[2].enq(req); //FIXME: replace with RXTX.
        end
      endcase
      // forward metadata to next stage.
      metadata_ff[1].enq(meta);
    end
  endrule

  rule rl_handle_response if (interruptStatus);
    let v <- toGet(bbRspFifo[readyChannel]).get;
    let meta <- toGet(metadata_ff[1]).get;
    case (v) matches
      tagged NopRspT {pkt: .pkt}: begin
        MetadataResponse rsp = tagged VlanDecapNopRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RemoveVlanSingleTaggedRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged VlanDecapRemoveVlanSingleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
      tagged RemoveVlanDoubleTaggedRspT {pkt: .pkt, ethernet$etherType: .ethernet$etherType}: begin
        meta.ethernet$etherType = tagged Valid ethernet$etherType;
        MetadataResponse rsp = tagged VlanDecapRemoveVlanDoubleTaggedRspT {pkt: pkt, meta: meta};
        tx_info_metadata.enq(rsp);
      end
    endcase
  endrule

  interface prev_control_state_0 = toServer(rx_metadata.e, tx_metadata.e);
  interface next_control_state_0 = toClient(bbReqFifo[0], bbRspFifo[0]);
  interface next_control_state_1 = toClient(bbReqFifo[1], bbRspFifo[1]);
  interface next_control_state_2 = toClient(bbReqFifo[2], bbRspFifo[2]);
endmodule

// ====== EGRESS ======

interface Egress;
  interface Client#(MetadataRequest, MetadataResponse) next;
endinterface
module mkEgress #(Vector#(numClients, Client#(MetadataRequest, MetadataResponse)) mdc) (Egress);
  FIFOF#(MetadataRequest) default_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) default_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) egress_acl_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) egress_acl_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) egress_bd_map_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) egress_bd_map_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) egress_bd_stats_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) egress_bd_stats_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) egress_filter_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) egress_filter_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) egress_filter_drop_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) egress_filter_drop_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) egress_port_mapping_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) egress_port_mapping_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) egress_vlan_xlate_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) egress_vlan_xlate_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) egress_vni_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) egress_vni_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_bos_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_bos_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_insert_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_insert_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_inst_0003_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_inst_0003_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_inst_0407_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_inst_0407_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_inst_0811_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_inst_0811_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_inst_1215_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_inst_1215_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_meta_header_update_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_meta_header_update_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) int_outer_encap_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) int_outer_encap_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) l3_rewrite_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) l3_rewrite_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) mirror_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) mirror_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) mtu_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) mtu_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) replica_type_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) replica_type_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) rewrite_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) rewrite_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) rewrite_multicast_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) rewrite_multicast_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) rid_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) rid_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) smac_rewrite_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) smac_rewrite_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_decap_process_inner_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_decap_process_inner_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_decap_process_outer_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_decap_process_outer_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_dmac_rewrite_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_dmac_rewrite_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_dst_rewrite_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_dst_rewrite_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_encap_process_inner_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_encap_process_inner_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_encap_process_outer_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_encap_process_outer_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_mtu_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_mtu_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_rewrite_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_rewrite_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_smac_rewrite_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_smac_rewrite_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) tunnel_src_rewrite_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) tunnel_src_rewrite_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) vlan_decap_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) vlan_decap_rsp_ff <- mkFIFOF;
  FIFOF#(MetadataRequest) next_req_ff <- mkFIFOF;
  FIFOF#(MetadataResponse) next_rsp_ff <- mkFIFOF;
  Vector#(numClients, Server#(MetadataRequest, MetadataResponse)) mds = replicate(toServer(default_req_ff, default_rsp_ff));
  mkConnection(mds, mdc);
  EgressAcl egress_acl <- mkEgressAcl();
  EgressBdMap egress_bd_map <- mkEgressBdMap();
  EgressBdStats egress_bd_stats <- mkEgressBdStats();
  EgressFilter egress_filter <- mkEgressFilter();
  EgressFilterDrop egress_filter_drop <- mkEgressFilterDrop();
  EgressPortMapping egress_port_mapping <- mkEgressPortMapping();
  EgressVlanXlate egress_vlan_xlate <- mkEgressVlanXlate();
  EgressVni egress_vni <- mkEgressVni();
  IntBos int_bos <- mkIntBos();
  IntInsert int_insert <- mkIntInsert();
  IntInst0003 int_inst_0003 <- mkIntInst0003();
  IntInst0407 int_inst_0407 <- mkIntInst0407();
  IntInst0811 int_inst_0811 <- mkIntInst0811();
  IntInst1215 int_inst_1215 <- mkIntInst1215();
  IntMetaHeaderUpdate int_meta_header_update <- mkIntMetaHeaderUpdate();
  IntOuterEncap int_outer_encap <- mkIntOuterEncap();
  L3Rewrite l3_rewrite <- mkL3Rewrite();
  Mirror mirror <- mkMirror();
  Mtu mtu <- mkMtu();
  ReplicaType replica_type <- mkReplicaType();
  Rewrite rewrite <- mkRewrite();
  RewriteMulticast rewrite_multicast <- mkRewriteMulticast();
  Rid rid <- mkRid();
  SmacRewrite smac_rewrite <- mkSmacRewrite();
  TunnelDecapProcessInner tunnel_decap_process_inner <- mkTunnelDecapProcessInner();
  TunnelDecapProcessOuter tunnel_decap_process_outer <- mkTunnelDecapProcessOuter();
  TunnelDmacRewrite tunnel_dmac_rewrite <- mkTunnelDmacRewrite();
  TunnelDstRewrite tunnel_dst_rewrite <- mkTunnelDstRewrite();
  TunnelEncapProcessInner tunnel_encap_process_inner <- mkTunnelEncapProcessInner();
  TunnelEncapProcessOuter tunnel_encap_process_outer <- mkTunnelEncapProcessOuter();
  TunnelMtu tunnel_mtu <- mkTunnelMtu();
  TunnelRewrite tunnel_rewrite <- mkTunnelRewrite();
  TunnelSmacRewrite tunnel_smac_rewrite <- mkTunnelSmacRewrite();
  TunnelSrcRewrite tunnel_src_rewrite <- mkTunnelSrcRewrite();
  VlanDecap vlan_decap <- mkVlanDecap();
  mkConnection(toClient(egress_acl_req_ff, egress_acl_rsp_ff), egress_acl.prev_control_state_0);
  mkConnection(toClient(egress_bd_map_req_ff, egress_bd_map_rsp_ff), egress_bd_map.prev_control_state_0);
  mkConnection(toClient(egress_bd_stats_req_ff, egress_bd_stats_rsp_ff), egress_bd_stats.prev_control_state_0);
  mkConnection(toClient(egress_filter_req_ff, egress_filter_rsp_ff), egress_filter.prev_control_state_0);
  mkConnection(toClient(egress_filter_drop_req_ff, egress_filter_drop_rsp_ff), egress_filter_drop.prev_control_state_0);
  mkConnection(toClient(egress_port_mapping_req_ff, egress_port_mapping_rsp_ff), egress_port_mapping.prev_control_state_0);
  mkConnection(toClient(egress_vlan_xlate_req_ff, egress_vlan_xlate_rsp_ff), egress_vlan_xlate.prev_control_state_0);
  mkConnection(toClient(egress_vni_req_ff, egress_vni_rsp_ff), egress_vni.prev_control_state_0);
  mkConnection(toClient(int_bos_req_ff, int_bos_rsp_ff), int_bos.prev_control_state_0);
  mkConnection(toClient(int_insert_req_ff, int_insert_rsp_ff), int_insert.prev_control_state_0);
  mkConnection(toClient(int_inst_0003_req_ff, int_inst_0003_rsp_ff), int_inst_0003.prev_control_state_0);
  mkConnection(toClient(int_inst_0407_req_ff, int_inst_0407_rsp_ff), int_inst_0407.prev_control_state_0);
  mkConnection(toClient(int_inst_0811_req_ff, int_inst_0811_rsp_ff), int_inst_0811.prev_control_state_0);
  mkConnection(toClient(int_inst_1215_req_ff, int_inst_1215_rsp_ff), int_inst_1215.prev_control_state_0);
  mkConnection(toClient(int_meta_header_update_req_ff, int_meta_header_update_rsp_ff), int_meta_header_update.prev_control_state_0);
  mkConnection(toClient(int_outer_encap_req_ff, int_outer_encap_rsp_ff), int_outer_encap.prev_control_state_0);
  mkConnection(toClient(l3_rewrite_req_ff, l3_rewrite_rsp_ff), l3_rewrite.prev_control_state_0);
  mkConnection(toClient(mirror_req_ff, mirror_rsp_ff), mirror.prev_control_state_0);
  mkConnection(toClient(mtu_req_ff, mtu_rsp_ff), mtu.prev_control_state_0);
  mkConnection(toClient(replica_type_req_ff, replica_type_rsp_ff), replica_type.prev_control_state_0);
  mkConnection(toClient(rewrite_req_ff, rewrite_rsp_ff), rewrite.prev_control_state_0);
  mkConnection(toClient(rewrite_multicast_req_ff, rewrite_multicast_rsp_ff), rewrite_multicast.prev_control_state_0);
  mkConnection(toClient(rid_req_ff, rid_rsp_ff), rid.prev_control_state_0);
  mkConnection(toClient(smac_rewrite_req_ff, smac_rewrite_rsp_ff), smac_rewrite.prev_control_state_0);
  mkConnection(toClient(tunnel_decap_process_inner_req_ff, tunnel_decap_process_inner_rsp_ff), tunnel_decap_process_inner.prev_control_state_0);
  mkConnection(toClient(tunnel_decap_process_outer_req_ff, tunnel_decap_process_outer_rsp_ff), tunnel_decap_process_outer.prev_control_state_0);
  mkConnection(toClient(tunnel_dmac_rewrite_req_ff, tunnel_dmac_rewrite_rsp_ff), tunnel_dmac_rewrite.prev_control_state_0);
  mkConnection(toClient(tunnel_dst_rewrite_req_ff, tunnel_dst_rewrite_rsp_ff), tunnel_dst_rewrite.prev_control_state_0);
  mkConnection(toClient(tunnel_encap_process_inner_req_ff, tunnel_encap_process_inner_rsp_ff), tunnel_encap_process_inner.prev_control_state_0);
  mkConnection(toClient(tunnel_encap_process_outer_req_ff, tunnel_encap_process_outer_rsp_ff), tunnel_encap_process_outer.prev_control_state_0);
  mkConnection(toClient(tunnel_mtu_req_ff, tunnel_mtu_rsp_ff), tunnel_mtu.prev_control_state_0);
  mkConnection(toClient(tunnel_rewrite_req_ff, tunnel_rewrite_rsp_ff), tunnel_rewrite.prev_control_state_0);
  mkConnection(toClient(tunnel_smac_rewrite_req_ff, tunnel_smac_rewrite_rsp_ff), tunnel_smac_rewrite.prev_control_state_0);
  mkConnection(toClient(tunnel_src_rewrite_req_ff, tunnel_src_rewrite_rsp_ff), tunnel_src_rewrite.prev_control_state_0);
  mkConnection(toClient(vlan_decap_req_ff, vlan_decap_rsp_ff), vlan_decap.prev_control_state_0);
  // Basic Blocks
  Nop nop_0 <- mkNop();
  EgressMirror egress_mirror_0 <- mkEgressMirror();
  EgressMirrorDrop egress_mirror_drop_0 <- mkEgressMirrorDrop();
  EgressRedirectToCpu egress_redirect_to_cpu_0 <- mkEgressRedirectToCpu();
  Nop nop_1 <- mkNop();
  SetEgressBdProperties set_egress_bd_properties_0 <- mkSetEgressBdProperties();
  Nop nop_2 <- mkNop();
  EgressFilterCheck egress_filter_check_0 <- mkEgressFilterCheck();
  SetEgressFilterDrop set_egress_filter_drop_0 <- mkSetEgressFilterDrop();
  EgressPortTypeNormal egress_port_type_normal_0 <- mkEgressPortTypeNormal();
  EgressPortTypeFabric egress_port_type_fabric_0 <- mkEgressPortTypeFabric();
  EgressPortTypeCpu egress_port_type_cpu_0 <- mkEgressPortTypeCpu();
  SetEgressPacketVlanUntagged set_egress_packet_vlan_untagged_0 <- mkSetEgressPacketVlanUntagged();
  SetEgressPacketVlanTagged set_egress_packet_vlan_tagged_0 <- mkSetEgressPacketVlanTagged();
  SetEgressPacketVlanDoubleTagged set_egress_packet_vlan_double_tagged_0 <- mkSetEgressPacketVlanDoubleTagged();
  Nop nop_3 <- mkNop();
  SetEgressTunnelVni set_egress_tunnel_vni_0 <- mkSetEgressTunnelVni();
  IntSetHeader0Bos int_set_header_0_bos_0 <- mkIntSetHeader0Bos();
  IntSetHeader1Bos int_set_header_1_bos_0 <- mkIntSetHeader1Bos();
  IntSetHeader2Bos int_set_header_2_bos_0 <- mkIntSetHeader2Bos();
  IntSetHeader3Bos int_set_header_3_bos_0 <- mkIntSetHeader3Bos();
  IntSetHeader4Bos int_set_header_4_bos_0 <- mkIntSetHeader4Bos();
  IntSetHeader5Bos int_set_header_5_bos_0 <- mkIntSetHeader5Bos();
  IntSetHeader6Bos int_set_header_6_bos_0 <- mkIntSetHeader6Bos();
  IntSetHeader7Bos int_set_header_7_bos_0 <- mkIntSetHeader7Bos();
  Nop nop_4 <- mkNop();
  IntTransit int_transit_0 <- mkIntTransit();
  IntSrc int_src_0 <- mkIntSrc();
  IntReset int_reset_0 <- mkIntReset();
  IntSetHeader0003I0 int_set_header_0003_i0_0 <- mkIntSetHeader0003I0();
  IntSetHeader0003I1 int_set_header_0003_i1_0 <- mkIntSetHeader0003I1();
  IntSetHeader0003I2 int_set_header_0003_i2_0 <- mkIntSetHeader0003I2();
  IntSetHeader0003I3 int_set_header_0003_i3_0 <- mkIntSetHeader0003I3();
  IntSetHeader0003I4 int_set_header_0003_i4_0 <- mkIntSetHeader0003I4();
  IntSetHeader0003I5 int_set_header_0003_i5_0 <- mkIntSetHeader0003I5();
  IntSetHeader0003I6 int_set_header_0003_i6_0 <- mkIntSetHeader0003I6();
  IntSetHeader0003I7 int_set_header_0003_i7_0 <- mkIntSetHeader0003I7();
  IntSetHeader0003I8 int_set_header_0003_i8_0 <- mkIntSetHeader0003I8();
  IntSetHeader0003I9 int_set_header_0003_i9_0 <- mkIntSetHeader0003I9();
  IntSetHeader0003I10 int_set_header_0003_i10_0 <- mkIntSetHeader0003I10();
  IntSetHeader0003I11 int_set_header_0003_i11_0 <- mkIntSetHeader0003I11();
  IntSetHeader0003I12 int_set_header_0003_i12_0 <- mkIntSetHeader0003I12();
  IntSetHeader0003I13 int_set_header_0003_i13_0 <- mkIntSetHeader0003I13();
  IntSetHeader0003I14 int_set_header_0003_i14_0 <- mkIntSetHeader0003I14();
  IntSetHeader0003I15 int_set_header_0003_i15_0 <- mkIntSetHeader0003I15();
  IntSetHeader0407I0 int_set_header_0407_i0_0 <- mkIntSetHeader0407I0();
  IntSetHeader0407I1 int_set_header_0407_i1_0 <- mkIntSetHeader0407I1();
  IntSetHeader0407I2 int_set_header_0407_i2_0 <- mkIntSetHeader0407I2();
  IntSetHeader0407I3 int_set_header_0407_i3_0 <- mkIntSetHeader0407I3();
  IntSetHeader0407I4 int_set_header_0407_i4_0 <- mkIntSetHeader0407I4();
  IntSetHeader0407I5 int_set_header_0407_i5_0 <- mkIntSetHeader0407I5();
  IntSetHeader0407I6 int_set_header_0407_i6_0 <- mkIntSetHeader0407I6();
  IntSetHeader0407I7 int_set_header_0407_i7_0 <- mkIntSetHeader0407I7();
  IntSetHeader0407I8 int_set_header_0407_i8_0 <- mkIntSetHeader0407I8();
  IntSetHeader0407I9 int_set_header_0407_i9_0 <- mkIntSetHeader0407I9();
  IntSetHeader0407I10 int_set_header_0407_i10_0 <- mkIntSetHeader0407I10();
  IntSetHeader0407I11 int_set_header_0407_i11_0 <- mkIntSetHeader0407I11();
  IntSetHeader0407I12 int_set_header_0407_i12_0 <- mkIntSetHeader0407I12();
  IntSetHeader0407I13 int_set_header_0407_i13_0 <- mkIntSetHeader0407I13();
  IntSetHeader0407I14 int_set_header_0407_i14_0 <- mkIntSetHeader0407I14();
  IntSetHeader0407I15 int_set_header_0407_i15_0 <- mkIntSetHeader0407I15();
  Nop nop_5 <- mkNop();
  Nop nop_6 <- mkNop();
  Nop nop_7 <- mkNop();
  IntSetEBit int_set_e_bit_0 <- mkIntSetEBit();
  IntUpdateTotalHopCnt int_update_total_hop_cnt_0 <- mkIntUpdateTotalHopCnt();
  IntUpdateVxlanGpeIpv4 int_update_vxlan_gpe_ipv4_0 <- mkIntUpdateVxlanGpeIpv4();
  IntAddUpdateVxlanGpeIpv4 int_add_update_vxlan_gpe_ipv4_0 <- mkIntAddUpdateVxlanGpeIpv4();
  Nop nop_8 <- mkNop();
  Nop nop_9 <- mkNop();
  Ipv4UnicastRewrite ipv4_unicast_rewrite_0 <- mkIpv4UnicastRewrite();
  Ipv4MulticastRewrite ipv4_multicast_rewrite_0 <- mkIpv4MulticastRewrite();
  Ipv6UnicastRewrite ipv6_unicast_rewrite_0 <- mkIpv6UnicastRewrite();
  Ipv6MulticastRewrite ipv6_multicast_rewrite_0 <- mkIpv6MulticastRewrite();
  MplsRewrite mpls_rewrite_0 <- mkMplsRewrite();
  Nop nop_10 <- mkNop();
  SetMirrorNhop set_mirror_nhop_0 <- mkSetMirrorNhop();
  SetMirrorBd set_mirror_bd_0 <- mkSetMirrorBd();
  SflowPktToCpu sflow_pkt_to_cpu_0 <- mkSflowPktToCpu();
  MtuMiss mtu_miss_0 <- mkMtuMiss();
  Ipv4MtuCheck ipv4_mtu_check_0 <- mkIpv4MtuCheck();
  Ipv6MtuCheck ipv6_mtu_check_0 <- mkIpv6MtuCheck();
  Nop nop_11 <- mkNop();
  SetReplicaCopyBridged set_replica_copy_bridged_0 <- mkSetReplicaCopyBridged();
  Nop nop_12 <- mkNop();
  SetL2Rewrite set_l2_rewrite_0 <- mkSetL2Rewrite();
  SetL2RewriteWithTunnel set_l2_rewrite_with_tunnel_0 <- mkSetL2RewriteWithTunnel();
  SetL3Rewrite set_l3_rewrite_0 <- mkSetL3Rewrite();
  SetL3RewriteWithTunnel set_l3_rewrite_with_tunnel_0 <- mkSetL3RewriteWithTunnel();
  SetMplsSwapPushRewriteL2 set_mpls_swap_push_rewrite_l2_0 <- mkSetMplsSwapPushRewriteL2();
  SetMplsPushRewriteL2 set_mpls_push_rewrite_l2_0 <- mkSetMplsPushRewriteL2();
  SetMplsSwapPushRewriteL3 set_mpls_swap_push_rewrite_l3_0 <- mkSetMplsSwapPushRewriteL3();
  SetMplsPushRewriteL3 set_mpls_push_rewrite_l3_0 <- mkSetMplsPushRewriteL3();
  Nop nop_13 <- mkNop();
  RewriteIpv4Multicast rewrite_ipv4_multicast_0 <- mkRewriteIpv4Multicast();
  RewriteIpv6Multicast rewrite_ipv6_multicast_0 <- mkRewriteIpv6Multicast();
  Nop nop_14 <- mkNop();
  OuterReplicaFromRid outer_replica_from_rid_0 <- mkOuterReplicaFromRid();
  InnerReplicaFromRid inner_replica_from_rid_0 <- mkInnerReplicaFromRid();
  RewriteSmac rewrite_smac_0 <- mkRewriteSmac();
  DecapInnerUdp decap_inner_udp_0 <- mkDecapInnerUdp();
  DecapInnerTcp decap_inner_tcp_0 <- mkDecapInnerTcp();
  DecapInnerIcmp decap_inner_icmp_0 <- mkDecapInnerIcmp();
  DecapInnerUnknown decap_inner_unknown_0 <- mkDecapInnerUnknown();
  DecapVxlanInnerIpv4 decap_vxlan_inner_ipv4_0 <- mkDecapVxlanInnerIpv4();
  DecapVxlanInnerIpv6 decap_vxlan_inner_ipv6_0 <- mkDecapVxlanInnerIpv6();
  DecapVxlanInnerNonIp decap_vxlan_inner_non_ip_0 <- mkDecapVxlanInnerNonIp();
  DecapGenvInnerIpv4 decap_genv_inner_ipv4_0 <- mkDecapGenvInnerIpv4();
  DecapGenvInnerIpv6 decap_genv_inner_ipv6_0 <- mkDecapGenvInnerIpv6();
  DecapGenvInnerNonIp decap_genv_inner_non_ip_0 <- mkDecapGenvInnerNonIp();
  DecapNvgreInnerIpv4 decap_nvgre_inner_ipv4_0 <- mkDecapNvgreInnerIpv4();
  DecapNvgreInnerIpv6 decap_nvgre_inner_ipv6_0 <- mkDecapNvgreInnerIpv6();
  DecapNvgreInnerNonIp decap_nvgre_inner_non_ip_0 <- mkDecapNvgreInnerNonIp();
  DecapGreInnerIpv4 decap_gre_inner_ipv4_0 <- mkDecapGreInnerIpv4();
  DecapGreInnerIpv6 decap_gre_inner_ipv6_0 <- mkDecapGreInnerIpv6();
  DecapGreInnerNonIp decap_gre_inner_non_ip_0 <- mkDecapGreInnerNonIp();
  DecapIpInnerIpv4 decap_ip_inner_ipv4_0 <- mkDecapIpInnerIpv4();
  DecapIpInnerIpv6 decap_ip_inner_ipv6_0 <- mkDecapIpInnerIpv6();
  DecapMplsInnerIpv4Pop1 decap_mpls_inner_ipv4_pop1_0 <- mkDecapMplsInnerIpv4Pop1();
  DecapMplsInnerIpv6Pop1 decap_mpls_inner_ipv6_pop1_0 <- mkDecapMplsInnerIpv6Pop1();
  DecapMplsInnerEthernetIpv4Pop1 decap_mpls_inner_ethernet_ipv4_pop1_0 <- mkDecapMplsInnerEthernetIpv4Pop1();
  DecapMplsInnerEthernetIpv6Pop1 decap_mpls_inner_ethernet_ipv6_pop1_0 <- mkDecapMplsInnerEthernetIpv6Pop1();
  DecapMplsInnerEthernetNonIpPop1 decap_mpls_inner_ethernet_non_ip_pop1_0 <- mkDecapMplsInnerEthernetNonIpPop1();
  DecapMplsInnerIpv4Pop2 decap_mpls_inner_ipv4_pop2_0 <- mkDecapMplsInnerIpv4Pop2();
  DecapMplsInnerIpv6Pop2 decap_mpls_inner_ipv6_pop2_0 <- mkDecapMplsInnerIpv6Pop2();
  DecapMplsInnerEthernetIpv4Pop2 decap_mpls_inner_ethernet_ipv4_pop2_0 <- mkDecapMplsInnerEthernetIpv4Pop2();
  DecapMplsInnerEthernetIpv6Pop2 decap_mpls_inner_ethernet_ipv6_pop2_0 <- mkDecapMplsInnerEthernetIpv6Pop2();
  DecapMplsInnerEthernetNonIpPop2 decap_mpls_inner_ethernet_non_ip_pop2_0 <- mkDecapMplsInnerEthernetNonIpPop2();
  DecapMplsInnerIpv4Pop3 decap_mpls_inner_ipv4_pop3_0 <- mkDecapMplsInnerIpv4Pop3();
  DecapMplsInnerIpv6Pop3 decap_mpls_inner_ipv6_pop3_0 <- mkDecapMplsInnerIpv6Pop3();
  DecapMplsInnerEthernetIpv4Pop3 decap_mpls_inner_ethernet_ipv4_pop3_0 <- mkDecapMplsInnerEthernetIpv4Pop3();
  DecapMplsInnerEthernetIpv6Pop3 decap_mpls_inner_ethernet_ipv6_pop3_0 <- mkDecapMplsInnerEthernetIpv6Pop3();
  DecapMplsInnerEthernetNonIpPop3 decap_mpls_inner_ethernet_non_ip_pop3_0 <- mkDecapMplsInnerEthernetNonIpPop3();
  Nop nop_15 <- mkNop();
  RewriteTunnelDmac rewrite_tunnel_dmac_0 <- mkRewriteTunnelDmac();
  Nop nop_16 <- mkNop();
  RewriteTunnelIpv4Dst rewrite_tunnel_ipv4_dst_0 <- mkRewriteTunnelIpv4Dst();
  RewriteTunnelIpv6Dst rewrite_tunnel_ipv6_dst_0 <- mkRewriteTunnelIpv6Dst();
  InnerIpv4UdpRewrite inner_ipv4_udp_rewrite_0 <- mkInnerIpv4UdpRewrite();
  InnerIpv4TcpRewrite inner_ipv4_tcp_rewrite_0 <- mkInnerIpv4TcpRewrite();
  InnerIpv4IcmpRewrite inner_ipv4_icmp_rewrite_0 <- mkInnerIpv4IcmpRewrite();
  InnerIpv4UnknownRewrite inner_ipv4_unknown_rewrite_0 <- mkInnerIpv4UnknownRewrite();
  InnerIpv6UdpRewrite inner_ipv6_udp_rewrite_0 <- mkInnerIpv6UdpRewrite();
  InnerIpv6TcpRewrite inner_ipv6_tcp_rewrite_0 <- mkInnerIpv6TcpRewrite();
  InnerIpv6IcmpRewrite inner_ipv6_icmp_rewrite_0 <- mkInnerIpv6IcmpRewrite();
  InnerIpv6UnknownRewrite inner_ipv6_unknown_rewrite_0 <- mkInnerIpv6UnknownRewrite();
  InnerNonIpRewrite inner_non_ip_rewrite_0 <- mkInnerNonIpRewrite();
  Nop nop_17 <- mkNop();
  Ipv4VxlanRewrite ipv4_vxlan_rewrite_0 <- mkIpv4VxlanRewrite();
  Ipv4GenvRewrite ipv4_genv_rewrite_0 <- mkIpv4GenvRewrite();
  Ipv4NvgreRewrite ipv4_nvgre_rewrite_0 <- mkIpv4NvgreRewrite();
  Ipv4GreRewrite ipv4_gre_rewrite_0 <- mkIpv4GreRewrite();
  Ipv4IpRewrite ipv4_ip_rewrite_0 <- mkIpv4IpRewrite();
  Ipv4ErspanT3Rewrite ipv4_erspan_t3_rewrite_0 <- mkIpv4ErspanT3Rewrite();
  Ipv6GreRewrite ipv6_gre_rewrite_0 <- mkIpv6GreRewrite();
  Ipv6IpRewrite ipv6_ip_rewrite_0 <- mkIpv6IpRewrite();
  Ipv6NvgreRewrite ipv6_nvgre_rewrite_0 <- mkIpv6NvgreRewrite();
  Ipv6VxlanRewrite ipv6_vxlan_rewrite_0 <- mkIpv6VxlanRewrite();
  Ipv6GenvRewrite ipv6_genv_rewrite_0 <- mkIpv6GenvRewrite();
  Ipv6ErspanT3Rewrite ipv6_erspan_t3_rewrite_0 <- mkIpv6ErspanT3Rewrite();
  MplsEthernetPush1Rewrite mpls_ethernet_push1_rewrite_0 <- mkMplsEthernetPush1Rewrite();
  MplsIpPush1Rewrite mpls_ip_push1_rewrite_0 <- mkMplsIpPush1Rewrite();
  MplsEthernetPush2Rewrite mpls_ethernet_push2_rewrite_0 <- mkMplsEthernetPush2Rewrite();
  MplsIpPush2Rewrite mpls_ip_push2_rewrite_0 <- mkMplsIpPush2Rewrite();
  MplsEthernetPush3Rewrite mpls_ethernet_push3_rewrite_0 <- mkMplsEthernetPush3Rewrite();
  MplsIpPush3Rewrite mpls_ip_push3_rewrite_0 <- mkMplsIpPush3Rewrite();
  FabricRewrite fabric_rewrite_0 <- mkFabricRewrite();
  TunnelMtuCheck tunnel_mtu_check_0 <- mkTunnelMtuCheck();
  TunnelMtuMiss tunnel_mtu_miss_0 <- mkTunnelMtuMiss();
  Nop nop_18 <- mkNop();
  SetTunnelRewriteDetails set_tunnel_rewrite_details_0 <- mkSetTunnelRewriteDetails();
  SetMplsRewritePush1 set_mpls_rewrite_push1_0 <- mkSetMplsRewritePush1();
  SetMplsRewritePush2 set_mpls_rewrite_push2_0 <- mkSetMplsRewritePush2();
  SetMplsRewritePush3 set_mpls_rewrite_push3_0 <- mkSetMplsRewritePush3();
  CpuRxRewrite cpu_rx_rewrite_0 <- mkCpuRxRewrite();
  FabricUnicastRewrite fabric_unicast_rewrite_0 <- mkFabricUnicastRewrite();
  FabricMulticastRewrite fabric_multicast_rewrite_0 <- mkFabricMulticastRewrite();
  Nop nop_19 <- mkNop();
  RewriteTunnelSmac rewrite_tunnel_smac_0 <- mkRewriteTunnelSmac();
  Nop nop_20 <- mkNop();
  RewriteTunnelIpv4Src rewrite_tunnel_ipv4_src_0 <- mkRewriteTunnelIpv4Src();
  RewriteTunnelIpv6Src rewrite_tunnel_ipv6_src_0 <- mkRewriteTunnelIpv6Src();
  Nop nop_21 <- mkNop();
  RemoveVlanSingleTagged remove_vlan_single_tagged_0 <- mkRemoveVlanSingleTagged();
  RemoveVlanDoubleTagged remove_vlan_double_tagged_0 <- mkRemoveVlanDoubleTagged();
  mkChan(mkFIFOF, mkFIFOF, egress_acl.next_control_state_0, nop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_acl.next_control_state_1, egress_mirror_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_acl.next_control_state_2, egress_mirror_drop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_acl.next_control_state_3, egress_redirect_to_cpu_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_bd_map.next_control_state_0, nop_1.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_bd_map.next_control_state_1, set_egress_bd_properties_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_bd_stats.next_control_state_0, nop_2.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_filter.next_control_state_0, egress_filter_check_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_filter_drop.next_control_state_0, set_egress_filter_drop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_port_mapping.next_control_state_0, egress_port_type_normal_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_port_mapping.next_control_state_1, egress_port_type_fabric_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_port_mapping.next_control_state_2, egress_port_type_cpu_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_vlan_xlate.next_control_state_0, set_egress_packet_vlan_untagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_vlan_xlate.next_control_state_1, set_egress_packet_vlan_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_vlan_xlate.next_control_state_2, set_egress_packet_vlan_double_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_vni.next_control_state_0, nop_3.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, egress_vni.next_control_state_1, set_egress_tunnel_vni_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_0, int_set_header_0_bos_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_1, int_set_header_1_bos_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_2, int_set_header_2_bos_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_3, int_set_header_3_bos_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_4, int_set_header_4_bos_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_5, int_set_header_5_bos_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_6, int_set_header_6_bos_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_7, int_set_header_7_bos_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_bos.next_control_state_8, nop_4.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_insert.next_control_state_0, int_transit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_insert.next_control_state_1, int_src_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_insert.next_control_state_2, int_reset_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_0, int_set_header_0003_i0_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_1, int_set_header_0003_i1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_2, int_set_header_0003_i2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_3, int_set_header_0003_i3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_4, int_set_header_0003_i4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_5, int_set_header_0003_i5_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_6, int_set_header_0003_i6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_7, int_set_header_0003_i7_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_8, int_set_header_0003_i8_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_9, int_set_header_0003_i9_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_10, int_set_header_0003_i10_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_11, int_set_header_0003_i11_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_12, int_set_header_0003_i12_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_13, int_set_header_0003_i13_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_14, int_set_header_0003_i14_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0003.next_control_state_15, int_set_header_0003_i15_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_0, int_set_header_0407_i0_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_1, int_set_header_0407_i1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_2, int_set_header_0407_i2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_3, int_set_header_0407_i3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_4, int_set_header_0407_i4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_5, int_set_header_0407_i5_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_6, int_set_header_0407_i6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_7, int_set_header_0407_i7_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_8, int_set_header_0407_i8_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_9, int_set_header_0407_i9_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_10, int_set_header_0407_i10_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_11, int_set_header_0407_i11_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_12, int_set_header_0407_i12_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_13, int_set_header_0407_i13_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_14, int_set_header_0407_i14_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_15, int_set_header_0407_i15_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0407.next_control_state_16, nop_5.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_0811.next_control_state_0, nop_6.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_inst_1215.next_control_state_0, nop_7.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_meta_header_update.next_control_state_0, int_set_e_bit_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_meta_header_update.next_control_state_1, int_update_total_hop_cnt_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_outer_encap.next_control_state_0, int_update_vxlan_gpe_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_outer_encap.next_control_state_1, int_add_update_vxlan_gpe_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, int_outer_encap.next_control_state_2, nop_8.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, l3_rewrite.next_control_state_0, nop_9.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, l3_rewrite.next_control_state_1, ipv4_unicast_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, l3_rewrite.next_control_state_2, ipv4_multicast_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, l3_rewrite.next_control_state_3, ipv6_unicast_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, l3_rewrite.next_control_state_4, ipv6_multicast_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, l3_rewrite.next_control_state_5, mpls_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mirror.next_control_state_0, nop_10.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mirror.next_control_state_1, set_mirror_nhop_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mirror.next_control_state_2, set_mirror_bd_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mirror.next_control_state_3, sflow_pkt_to_cpu_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mtu.next_control_state_0, mtu_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mtu.next_control_state_1, ipv4_mtu_check_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, mtu.next_control_state_2, ipv6_mtu_check_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, replica_type.next_control_state_0, nop_11.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, replica_type.next_control_state_1, set_replica_copy_bridged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_0, nop_12.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_1, set_l2_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_2, set_l2_rewrite_with_tunnel_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_3, set_l3_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_4, set_l3_rewrite_with_tunnel_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_5, set_mpls_swap_push_rewrite_l2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_6, set_mpls_push_rewrite_l2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_7, set_mpls_swap_push_rewrite_l3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite.next_control_state_8, set_mpls_push_rewrite_l3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite_multicast.next_control_state_0, nop_13.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite_multicast.next_control_state_1, rewrite_ipv4_multicast_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rewrite_multicast.next_control_state_2, rewrite_ipv6_multicast_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rid.next_control_state_0, nop_14.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rid.next_control_state_1, outer_replica_from_rid_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, rid.next_control_state_2, inner_replica_from_rid_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, smac_rewrite.next_control_state_0, rewrite_smac_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_inner.next_control_state_0, decap_inner_udp_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_inner.next_control_state_1, decap_inner_tcp_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_inner.next_control_state_2, decap_inner_icmp_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_inner.next_control_state_3, decap_inner_unknown_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_0, decap_vxlan_inner_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_1, decap_vxlan_inner_ipv6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_2, decap_vxlan_inner_non_ip_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_3, decap_genv_inner_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_4, decap_genv_inner_ipv6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_5, decap_genv_inner_non_ip_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_6, decap_nvgre_inner_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_7, decap_nvgre_inner_ipv6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_8, decap_nvgre_inner_non_ip_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_9, decap_gre_inner_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_10, decap_gre_inner_ipv6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_11, decap_gre_inner_non_ip_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_12, decap_ip_inner_ipv4_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_13, decap_ip_inner_ipv6_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_14, decap_mpls_inner_ipv4_pop1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_15, decap_mpls_inner_ipv6_pop1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_16, decap_mpls_inner_ethernet_ipv4_pop1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_17, decap_mpls_inner_ethernet_ipv6_pop1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_18, decap_mpls_inner_ethernet_non_ip_pop1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_19, decap_mpls_inner_ipv4_pop2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_20, decap_mpls_inner_ipv6_pop2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_21, decap_mpls_inner_ethernet_ipv4_pop2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_22, decap_mpls_inner_ethernet_ipv6_pop2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_23, decap_mpls_inner_ethernet_non_ip_pop2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_24, decap_mpls_inner_ipv4_pop3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_25, decap_mpls_inner_ipv6_pop3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_26, decap_mpls_inner_ethernet_ipv4_pop3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_27, decap_mpls_inner_ethernet_ipv6_pop3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_decap_process_outer.next_control_state_28, decap_mpls_inner_ethernet_non_ip_pop3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_dmac_rewrite.next_control_state_0, nop_15.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_dmac_rewrite.next_control_state_1, rewrite_tunnel_dmac_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_dst_rewrite.next_control_state_0, nop_16.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_dst_rewrite.next_control_state_1, rewrite_tunnel_ipv4_dst_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_dst_rewrite.next_control_state_2, rewrite_tunnel_ipv6_dst_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_0, inner_ipv4_udp_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_1, inner_ipv4_tcp_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_2, inner_ipv4_icmp_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_3, inner_ipv4_unknown_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_4, inner_ipv6_udp_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_5, inner_ipv6_tcp_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_6, inner_ipv6_icmp_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_7, inner_ipv6_unknown_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_inner.next_control_state_8, inner_non_ip_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_0, nop_17.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_1, ipv4_vxlan_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_2, ipv4_genv_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_3, ipv4_nvgre_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_4, ipv4_gre_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_5, ipv4_ip_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_6, ipv4_erspan_t3_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_7, ipv6_gre_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_8, ipv6_ip_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_9, ipv6_nvgre_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_10, ipv6_vxlan_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_11, ipv6_genv_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_12, ipv6_erspan_t3_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_13, mpls_ethernet_push1_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_14, mpls_ip_push1_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_15, mpls_ethernet_push2_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_16, mpls_ip_push2_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_17, mpls_ethernet_push3_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_18, mpls_ip_push3_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_encap_process_outer.next_control_state_19, fabric_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_mtu.next_control_state_0, tunnel_mtu_check_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_mtu.next_control_state_1, tunnel_mtu_miss_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_rewrite.next_control_state_0, nop_18.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_rewrite.next_control_state_1, set_tunnel_rewrite_details_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_rewrite.next_control_state_2, set_mpls_rewrite_push1_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_rewrite.next_control_state_3, set_mpls_rewrite_push2_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_rewrite.next_control_state_4, set_mpls_rewrite_push3_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_rewrite.next_control_state_5, cpu_rx_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_rewrite.next_control_state_6, fabric_unicast_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_rewrite.next_control_state_7, fabric_multicast_rewrite_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_smac_rewrite.next_control_state_0, nop_19.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_smac_rewrite.next_control_state_1, rewrite_tunnel_smac_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_src_rewrite.next_control_state_0, nop_20.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_src_rewrite.next_control_state_1, rewrite_tunnel_ipv4_src_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, tunnel_src_rewrite.next_control_state_2, rewrite_tunnel_ipv6_src_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, vlan_decap.next_control_state_0, nop_21.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, vlan_decap.next_control_state_1, remove_vlan_single_tagged_0.prev_control_state);
  mkChan(mkFIFOF, mkFIFOF, vlan_decap.next_control_state_2, remove_vlan_double_tagged_0.prev_control_state);
  rule default_next_state if (default_req_ff.notEmpty);
    default_req_ff.deq;
    let _req = default_req_ff.first;
    let meta = _req.meta;
    let pkt = _req.pkt;
    if (( ( intrinsic_metadata$deflection_flag == 'h0 ) && ( egress_metadata$bypass == 'h0 ) )) begin
      if (( ( standard_metadata$instance_type != 'h0 ) && ( standard_metadata$instance_type != 'h5 ) )) begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        mirror_req_ff.enq(req);
      end
      else begin
        if (( intrinsic_metadata$egress_rid != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rid_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_port_mapping_req_ff.enq(req);
        end
      end
    end
    else begin
      if (( egress_metadata$bypass == 'h0 )) begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_acl_req_ff.enq(req);
      end
    end
  endrule

  rule egress_acl_next_state if (egress_acl_rsp_ff.notEmpty);
    egress_acl_rsp_ff.deq;
    let _rsp = egress_acl_rsp_ff.first;
    case (_rsp) matches
      tagged EgressAclNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        next_req_ff.enq(req);
      end
      tagged EgressAclEgressMirrorRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        next_req_ff.enq(req);
      end
      tagged EgressAclEgressMirrorDropRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        next_req_ff.enq(req);
      end
      tagged EgressAclEgressRedirectToCpuRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        next_req_ff.enq(req);
      end
    endcase
  endrule

  rule egress_bd_map_next_state if (egress_bd_map_rsp_ff.notEmpty);
    egress_bd_map_rsp_ff.deq;
    let _rsp = egress_bd_map_rsp_ff.first;
    case (_rsp) matches
      tagged EgressBdMapNopRspT {meta: .meta, pkt: .pkt}: begin
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( egress_metadata$routed == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          l3_rewrite_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          mtu_req_ff.enq(req);
        end
      end
      tagged EgressBdMapSetEgressBdPropertiesRspT {meta: .meta, pkt: .pkt}: begin
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( egress_metadata$routed == 'h1 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          l3_rewrite_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          mtu_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule egress_bd_stats_next_state if (egress_bd_stats_rsp_ff.notEmpty);
    egress_bd_stats_rsp_ff.deq;
    let _rsp = egress_bd_stats_rsp_ff.first;
    case (_rsp) matches
      tagged EgressBdStatsNopRspT {meta: .meta, pkt: .pkt}: begin
        let int_metadata$insert_cnt = fromMaybe(?, meta.int_metadata$insert_cnt);
        let fabric_metadata$fabric_header_present = fromMaybe(?, meta.fabric_metadata$fabric_header_present);
        let egress_metadata$port_type = fromMaybe(?, meta.egress_metadata$port_type);
        let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
        if (( ( fabric_metadata$fabric_header_present == 'h0 ) && ( tunnel_metadata$egress_tunnel_type != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_vni_req_ff.enq(req);
        end
        else begin
          if (( int_metadata$insert_cnt != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            int_outer_encap_req_ff.enq(req);
          end
          else begin
            if (( egress_metadata$port_type == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              egress_vlan_xlate_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              egress_filter_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule egress_filter_next_state if (egress_filter_rsp_ff.notEmpty);
    egress_filter_rsp_ff.deq;
    let _rsp = egress_filter_rsp_ff.first;
    case (_rsp) matches
      tagged EgressFilterEgressFilterCheckRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
        let multicast_metadata$inner_replica = fromMaybe(?, meta.multicast_metadata$inner_replica);
        let tunnel_metadata$ingress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$ingress_tunnel_type);
        let egress_filter_metadata$inner_bd = fromMaybe(?, meta.egress_filter_metadata$inner_bd);
        let egress_metadata$bypass = fromMaybe(?, meta.egress_metadata$bypass);
        let egress_filter_metadata$bd = fromMaybe(?, meta.egress_filter_metadata$bd);
        let egress_filter_metadata$ifindex_check = fromMaybe(?, meta.egress_filter_metadata$ifindex_check);
        if (( multicast_metadata$inner_replica == 'h1 )) begin
          if (( ( ( ( ( tunnel_metadata$ingress_tunnel_type == 'h0 ) && ( tunnel_metadata$egress_tunnel_type == 'h0 ) ) && ( egress_filter_metadata$bd == 'h0 ) ) && ( egress_filter_metadata$ifindex_check == 'h0 ) ) || ( ( ( tunnel_metadata$ingress_tunnel_type != 'h0 ) && ( tunnel_metadata$egress_tunnel_type != 'h0 ) ) && ( egress_filter_metadata$inner_bd == 'h0 ) ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            egress_filter_drop_req_ff.enq(req);
          end
          else begin
            if (( egress_metadata$bypass == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              egress_acl_req_ff.enq(req);
            end
          end
        end
        else begin
          if (( egress_metadata$bypass == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            egress_acl_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule egress_filter_drop_next_state if (egress_filter_drop_rsp_ff.notEmpty);
    egress_filter_drop_rsp_ff.deq;
    let _rsp = egress_filter_drop_rsp_ff.first;
    case (_rsp) matches
      tagged EgressFilterDropSetEgressFilterDropRspT {meta: .meta, pkt: .pkt}: begin
        let egress_metadata$bypass = fromMaybe(?, meta.egress_metadata$bypass);
        if (( egress_metadata$bypass == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_acl_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule egress_port_mapping_next_state if (egress_port_mapping_rsp_ff.notEmpty);
    egress_port_mapping_rsp_ff.deq;
    let _rsp = egress_port_mapping_rsp_ff.first;
    case (_rsp) matches
      tagged EgressPortMappingEgressPortTypeNormalRspT {meta: .meta, pkt: .pkt}: begin
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
        let multicast_metadata$replica = fromMaybe(?, meta.multicast_metadata$replica);
        let multicast_metadata$inner_replica = fromMaybe(?, meta.multicast_metadata$inner_replica);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let standard_metadata$instance_type = fromMaybe(?, meta.standard_metadata$instance_type);
        if (( ( standard_metadata$instance_type == 'h0 ) || ( standard_metadata$instance_type == 'h5 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          vlan_decap_req_ff.enq(req);
        end
        else begin
          if (( tunnel_metadata$tunnel_terminate == 'h1 )) begin
            if (( ( multicast_metadata$inner_replica == 'h1 ) || ( multicast_metadata$replica == 'h0 ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              tunnel_decap_process_outer_req_ff.enq(req);
            end
            else begin
              if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                rewrite_req_ff.enq(req);
              end
              else begin
                MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
                rewrite_multicast_req_ff.enq(req);
              end
            end
          end
          else begin
            if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              rewrite_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              rewrite_multicast_req_ff.enq(req);
            end
          end
        end
      end
      tagged EgressPortMappingEgressPortTypeFabricRspT {meta: .meta, pkt: .pkt}: begin
        let int_metadata$insert_cnt = fromMaybe(?, meta.int_metadata$insert_cnt);
        let fabric_metadata$fabric_header_present = fromMaybe(?, meta.fabric_metadata$fabric_header_present);
        let egress_metadata$port_type = fromMaybe(?, meta.egress_metadata$port_type);
        let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
        if (( ( fabric_metadata$fabric_header_present == 'h0 ) && ( tunnel_metadata$egress_tunnel_type != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_vni_req_ff.enq(req);
        end
        else begin
          if (( int_metadata$insert_cnt != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            int_outer_encap_req_ff.enq(req);
          end
          else begin
            if (( egress_metadata$port_type == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              egress_vlan_xlate_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              egress_filter_req_ff.enq(req);
            end
          end
        end
      end
      tagged EgressPortMappingEgressPortTypeCpuRspT {meta: .meta, pkt: .pkt}: begin
        let int_metadata$insert_cnt = fromMaybe(?, meta.int_metadata$insert_cnt);
        let fabric_metadata$fabric_header_present = fromMaybe(?, meta.fabric_metadata$fabric_header_present);
        let egress_metadata$port_type = fromMaybe(?, meta.egress_metadata$port_type);
        let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
        if (( ( fabric_metadata$fabric_header_present == 'h0 ) && ( tunnel_metadata$egress_tunnel_type != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_vni_req_ff.enq(req);
        end
        else begin
          if (( int_metadata$insert_cnt != 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            int_outer_encap_req_ff.enq(req);
          end
          else begin
            if (( egress_metadata$port_type == 'h0 )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              egress_vlan_xlate_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              egress_filter_req_ff.enq(req);
            end
          end
        end
      end
    endcase
  endrule

  rule egress_vlan_xlate_next_state if (egress_vlan_xlate_rsp_ff.notEmpty);
    egress_vlan_xlate_rsp_ff.deq;
    let _rsp = egress_vlan_xlate_rsp_ff.first;
    case (_rsp) matches
      tagged EgressVlanXlateSetEgressPacketVlanUntaggedRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_filter_req_ff.enq(req);
      end
      tagged EgressVlanXlateSetEgressPacketVlanTaggedRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_filter_req_ff.enq(req);
      end
      tagged EgressVlanXlateSetEgressPacketVlanDoubleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_filter_req_ff.enq(req);
      end
    endcase
  endrule

  rule egress_vni_next_state if (egress_vni_rsp_ff.notEmpty);
    egress_vni_rsp_ff.deq;
    let _rsp = egress_vni_rsp_ff.first;
    case (_rsp) matches
      tagged EgressVniNopRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
        if (( ( tunnel_metadata$egress_tunnel_type != 'hf ) && ( tunnel_metadata$egress_tunnel_type != 'h10 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_encap_process_inner_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_encap_process_outer_req_ff.enq(req);
        end
      end
      tagged EgressVniSetEgressTunnelVniRspT {meta: .meta, pkt: .pkt}: begin
        let tunnel_metadata$egress_tunnel_type = fromMaybe(?, meta.tunnel_metadata$egress_tunnel_type);
        if (( ( tunnel_metadata$egress_tunnel_type != 'hf ) && ( tunnel_metadata$egress_tunnel_type != 'h10 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_encap_process_inner_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          tunnel_encap_process_outer_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule int_bos_next_state if (int_bos_rsp_ff.notEmpty);
    int_bos_rsp_ff.deq;
    let _rsp = int_bos_rsp_ff.first;
    case (_rsp) matches
      tagged IntBosIntSetHeader0BosRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
      tagged IntBosIntSetHeader1BosRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
      tagged IntBosIntSetHeader2BosRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
      tagged IntBosIntSetHeader3BosRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
      tagged IntBosIntSetHeader4BosRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
      tagged IntBosIntSetHeader5BosRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
      tagged IntBosIntSetHeader6BosRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
      tagged IntBosIntSetHeader7BosRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
      tagged IntBosNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_meta_header_update_req_ff.enq(req);
      end
    endcase
  endrule

  rule int_insert_next_state if (int_insert_rsp_ff.notEmpty);
    int_insert_rsp_ff.deq;
    let _rsp = int_insert_rsp_ff.first;
    case (_rsp) matches
      tagged IntInsertIntTransitRspT {meta: .meta, pkt: .pkt}: begin
        let int_metadata$insert_cnt = fromMaybe(?, meta.int_metadata$insert_cnt);
        if (( int_metadata$insert_cnt != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          int_inst_0003_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          int_meta_header_update_req_ff.enq(req);
        end
      end
      tagged IntInsertIntSrcRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_stats_req_ff.enq(req);
      end
      tagged IntInsertIntResetRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_stats_req_ff.enq(req);
      end
    endcase
  endrule

  rule int_inst_0003_next_state if (int_inst_0003_rsp_ff.notEmpty);
    int_inst_0003_rsp_ff.deq;
    let _rsp = int_inst_0003_rsp_ff.first;
    case (_rsp) matches
      tagged IntInst0003IntSetHeader0003I0RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I5RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I7RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I8RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I9RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I10RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I11RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I12RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I13RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I14RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
      tagged IntInst0003IntSetHeader0003I15RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0407_req_ff.enq(req);
      end
    endcase
  endrule

  rule int_inst_0407_next_state if (int_inst_0407_rsp_ff.notEmpty);
    int_inst_0407_rsp_ff.deq;
    let _rsp = int_inst_0407_rsp_ff.first;
    case (_rsp) matches
      tagged IntInst0407IntSetHeader0407I0RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I5RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I7RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I8RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I9RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I10RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I11RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I12RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I13RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I14RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407IntSetHeader0407I15RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
      tagged IntInst0407NopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_0811_req_ff.enq(req);
      end
    endcase
  endrule

  rule int_inst_0811_next_state if (int_inst_0811_rsp_ff.notEmpty);
    int_inst_0811_rsp_ff.deq;
    let _rsp = int_inst_0811_rsp_ff.first;
    case (_rsp) matches
      tagged IntInst0811NopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_inst_1215_req_ff.enq(req);
      end
    endcase
  endrule

  rule int_inst_1215_next_state if (int_inst_1215_rsp_ff.notEmpty);
    int_inst_1215_rsp_ff.deq;
    let _rsp = int_inst_1215_rsp_ff.first;
    case (_rsp) matches
      tagged IntInst1215NopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_bos_req_ff.enq(req);
      end
    endcase
  endrule

  rule int_meta_header_update_next_state if (int_meta_header_update_rsp_ff.notEmpty);
    int_meta_header_update_rsp_ff.deq;
    let _rsp = int_meta_header_update_rsp_ff.first;
    case (_rsp) matches
      tagged IntMetaHeaderUpdateIntSetEBitRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_stats_req_ff.enq(req);
      end
      tagged IntMetaHeaderUpdateIntUpdateTotalHopCntRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_stats_req_ff.enq(req);
      end
    endcase
  endrule

  rule int_outer_encap_next_state if (int_outer_encap_rsp_ff.notEmpty);
    int_outer_encap_rsp_ff.deq;
    let _rsp = int_outer_encap_rsp_ff.first;
    case (_rsp) matches
      tagged IntOuterEncapIntUpdateVxlanGpeIpv4RspT {meta: .meta, pkt: .pkt}: begin
        let egress_metadata$port_type = fromMaybe(?, meta.egress_metadata$port_type);
        if (( egress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_vlan_xlate_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_filter_req_ff.enq(req);
        end
      end
      tagged IntOuterEncapIntAddUpdateVxlanGpeIpv4RspT {meta: .meta, pkt: .pkt}: begin
        let egress_metadata$port_type = fromMaybe(?, meta.egress_metadata$port_type);
        if (( egress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_vlan_xlate_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_filter_req_ff.enq(req);
        end
      end
      tagged IntOuterEncapNopRspT {meta: .meta, pkt: .pkt}: begin
        let egress_metadata$port_type = fromMaybe(?, meta.egress_metadata$port_type);
        if (( egress_metadata$port_type == 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_vlan_xlate_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          egress_filter_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule l3_rewrite_next_state if (l3_rewrite_rsp_ff.notEmpty);
    l3_rewrite_rsp_ff.deq;
    let _rsp = l3_rewrite_rsp_ff.first;
    case (_rsp) matches
      tagged L3RewriteNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        smac_rewrite_req_ff.enq(req);
      end
      tagged L3RewriteIpv4UnicastRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        smac_rewrite_req_ff.enq(req);
      end
      tagged L3RewriteIpv4MulticastRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        smac_rewrite_req_ff.enq(req);
      end
      tagged L3RewriteIpv6UnicastRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        smac_rewrite_req_ff.enq(req);
      end
      tagged L3RewriteIpv6MulticastRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        smac_rewrite_req_ff.enq(req);
      end
      tagged L3RewriteMplsRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        smac_rewrite_req_ff.enq(req);
      end
    endcase
  endrule

  rule mirror_next_state if (mirror_rsp_ff.notEmpty);
    mirror_rsp_ff.deq;
    let _rsp = mirror_rsp_ff.first;
    case (_rsp) matches
      tagged MirrorNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_port_mapping_req_ff.enq(req);
      end
      tagged MirrorSetMirrorNhopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_port_mapping_req_ff.enq(req);
      end
      tagged MirrorSetMirrorBdRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_port_mapping_req_ff.enq(req);
      end
      tagged MirrorSflowPktToCpuRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_port_mapping_req_ff.enq(req);
      end
    endcase
  endrule

  rule mtu_next_state if (mtu_rsp_ff.notEmpty);
    mtu_rsp_ff.deq;
    let _rsp = mtu_rsp_ff.first;
    case (_rsp) matches
      tagged MtuMtuMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_insert_req_ff.enq(req);
      end
      tagged MtuIpv4MtuCheckRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_insert_req_ff.enq(req);
      end
      tagged MtuIpv6MtuCheckRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        int_insert_req_ff.enq(req);
      end
    endcase
  endrule

  rule replica_type_next_state if (replica_type_rsp_ff.notEmpty);
    replica_type_rsp_ff.deq;
    let _rsp = replica_type_rsp_ff.first;
    case (_rsp) matches
      tagged ReplicaTypeNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_port_mapping_req_ff.enq(req);
      end
      tagged ReplicaTypeSetReplicaCopyBridgedRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_port_mapping_req_ff.enq(req);
      end
    endcase
  endrule

  rule rewrite_next_state if (rewrite_rsp_ff.notEmpty);
    rewrite_rsp_ff.deq;
    let _rsp = rewrite_rsp_ff.first;
    case (_rsp) matches
      tagged RewriteNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteSetL2RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteSetL2RewriteWithTunnelRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteSetL3RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteSetL3RewriteWithTunnelRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteSetMplsSwapPushRewriteL2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteSetMplsPushRewriteL2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteSetMplsSwapPushRewriteL3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteSetMplsPushRewriteL3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
    endcase
  endrule

  rule rewrite_multicast_next_state if (rewrite_multicast_rsp_ff.notEmpty);
    rewrite_multicast_rsp_ff.deq;
    let _rsp = rewrite_multicast_rsp_ff.first;
    case (_rsp) matches
      tagged RewriteMulticastNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteMulticastRewriteIpv4MulticastRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
      tagged RewriteMulticastRewriteIpv6MulticastRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        egress_bd_map_req_ff.enq(req);
      end
    endcase
  endrule

  rule rid_next_state if (rid_rsp_ff.notEmpty);
    rid_rsp_ff.deq;
    let _rsp = rid_rsp_ff.first;
    case (_rsp) matches
      tagged RidNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        replica_type_req_ff.enq(req);
      end
      tagged RidOuterReplicaFromRidRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        replica_type_req_ff.enq(req);
      end
      tagged RidInnerReplicaFromRidRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        replica_type_req_ff.enq(req);
      end
    endcase
  endrule

  rule smac_rewrite_next_state if (smac_rewrite_rsp_ff.notEmpty);
    smac_rewrite_rsp_ff.deq;
    let _rsp = smac_rewrite_rsp_ff.first;
    case (_rsp) matches
      tagged SmacRewriteRewriteSmacRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        mtu_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_decap_process_inner_next_state if (tunnel_decap_process_inner_rsp_ff.notEmpty);
    tunnel_decap_process_inner_rsp_ff.deq;
    let _rsp = tunnel_decap_process_inner_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelDecapProcessInnerDecapInnerUdpRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rewrite_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rewrite_multicast_req_ff.enq(req);
        end
      end
      tagged TunnelDecapProcessInnerDecapInnerTcpRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rewrite_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rewrite_multicast_req_ff.enq(req);
        end
      end
      tagged TunnelDecapProcessInnerDecapInnerIcmpRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rewrite_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rewrite_multicast_req_ff.enq(req);
        end
      end
      tagged TunnelDecapProcessInnerDecapInnerUnknownRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rewrite_req_ff.enq(req);
        end
        else begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          rewrite_multicast_req_ff.enq(req);
        end
      end
    endcase
  endrule

  rule tunnel_decap_process_outer_next_state if (tunnel_decap_process_outer_rsp_ff.notEmpty);
    tunnel_decap_process_outer_rsp_ff.deq;
    let _rsp = tunnel_decap_process_outer_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelDecapProcessOuterDecapVxlanInnerIpv4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapVxlanInnerIpv6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapVxlanInnerNonIpRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapGenvInnerIpv4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapGenvInnerIpv6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapGenvInnerNonIpRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapNvgreInnerIpv4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapNvgreInnerIpv6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapNvgreInnerNonIpRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapGreInnerIpv4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapGreInnerIpv6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapGreInnerNonIpRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapIpInnerIpv4RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapIpInnerIpv6RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerIpv4Pop1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerIpv6Pop1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv4Pop1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv6Pop1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetNonIpPop1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerIpv4Pop2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerIpv6Pop2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv4Pop2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv6Pop2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetNonIpPop2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerIpv4Pop3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerIpv6Pop3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv4Pop3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetIpv6Pop3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
      tagged TunnelDecapProcessOuterDecapMplsInnerEthernetNonIpPop3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_decap_process_inner_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_dmac_rewrite_next_state if (tunnel_dmac_rewrite_rsp_ff.notEmpty);
    tunnel_dmac_rewrite_rsp_ff.deq;
    let _rsp = tunnel_dmac_rewrite_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelDmacRewriteNopRspT {meta: .meta, pkt: .pkt}: begin
        let int_metadata$insert_cnt = fromMaybe(?, meta.int_metadata$insert_cnt);
        let egress_metadata$port_type = fromMaybe(?, meta.egress_metadata$port_type);
        if (( int_metadata$insert_cnt != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          int_outer_encap_req_ff.enq(req);
        end
        else begin
          if (( egress_metadata$port_type == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            egress_vlan_xlate_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            egress_filter_req_ff.enq(req);
          end
        end
      end
      tagged TunnelDmacRewriteRewriteTunnelDmacRspT {meta: .meta, pkt: .pkt}: begin
        let int_metadata$insert_cnt = fromMaybe(?, meta.int_metadata$insert_cnt);
        let egress_metadata$port_type = fromMaybe(?, meta.egress_metadata$port_type);
        if (( int_metadata$insert_cnt != 'h0 )) begin
          MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
          int_outer_encap_req_ff.enq(req);
        end
        else begin
          if (( egress_metadata$port_type == 'h0 )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            egress_vlan_xlate_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            egress_filter_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  rule tunnel_dst_rewrite_next_state if (tunnel_dst_rewrite_rsp_ff.notEmpty);
    tunnel_dst_rewrite_rsp_ff.deq;
    let _rsp = tunnel_dst_rewrite_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelDstRewriteNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_smac_rewrite_req_ff.enq(req);
      end
      tagged TunnelDstRewriteRewriteTunnelIpv4DstRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_smac_rewrite_req_ff.enq(req);
      end
      tagged TunnelDstRewriteRewriteTunnelIpv6DstRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_smac_rewrite_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_encap_process_inner_next_state if (tunnel_encap_process_inner_rsp_ff.notEmpty);
    tunnel_encap_process_inner_rsp_ff.deq;
    let _rsp = tunnel_encap_process_inner_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelEncapProcessInnerInnerIpv4UdpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
      tagged TunnelEncapProcessInnerInnerIpv4TcpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
      tagged TunnelEncapProcessInnerInnerIpv4IcmpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
      tagged TunnelEncapProcessInnerInnerIpv4UnknownRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
      tagged TunnelEncapProcessInnerInnerIpv6UdpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
      tagged TunnelEncapProcessInnerInnerIpv6TcpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
      tagged TunnelEncapProcessInnerInnerIpv6IcmpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
      tagged TunnelEncapProcessInnerInnerIpv6UnknownRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
      tagged TunnelEncapProcessInnerInnerNonIpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_encap_process_outer_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_encap_process_outer_next_state if (tunnel_encap_process_outer_rsp_ff.notEmpty);
    tunnel_encap_process_outer_rsp_ff.deq;
    let _rsp = tunnel_encap_process_outer_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelEncapProcessOuterNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv4VxlanRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv4GenvRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv4NvgreRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv4GreRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv4IpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv4ErspanT3RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv6GreRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv6IpRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv6NvgreRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv6VxlanRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv6GenvRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterIpv6ErspanT3RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterMplsEthernetPush1RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterMplsIpPush1RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterMplsEthernetPush2RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterMplsIpPush2RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterMplsEthernetPush3RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterMplsIpPush3RewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
      tagged TunnelEncapProcessOuterFabricRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_rewrite_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_mtu_next_state if (tunnel_mtu_rsp_ff.notEmpty);
    tunnel_mtu_rsp_ff.deq;
    let _rsp = tunnel_mtu_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelMtuTunnelMtuCheckRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_src_rewrite_req_ff.enq(req);
      end
      tagged TunnelMtuTunnelMtuMissRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_src_rewrite_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_rewrite_next_state if (tunnel_rewrite_rsp_ff.notEmpty);
    tunnel_rewrite_rsp_ff.deq;
    let _rsp = tunnel_rewrite_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelRewriteNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_mtu_req_ff.enq(req);
      end
      tagged TunnelRewriteSetTunnelRewriteDetailsRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_mtu_req_ff.enq(req);
      end
      tagged TunnelRewriteSetMplsRewritePush1RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_mtu_req_ff.enq(req);
      end
      tagged TunnelRewriteSetMplsRewritePush2RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_mtu_req_ff.enq(req);
      end
      tagged TunnelRewriteSetMplsRewritePush3RspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_mtu_req_ff.enq(req);
      end
      tagged TunnelRewriteCpuRxRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_mtu_req_ff.enq(req);
      end
      tagged TunnelRewriteFabricUnicastRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_mtu_req_ff.enq(req);
      end
      tagged TunnelRewriteFabricMulticastRewriteRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_mtu_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_smac_rewrite_next_state if (tunnel_smac_rewrite_rsp_ff.notEmpty);
    tunnel_smac_rewrite_rsp_ff.deq;
    let _rsp = tunnel_smac_rewrite_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelSmacRewriteNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_dmac_rewrite_req_ff.enq(req);
      end
      tagged TunnelSmacRewriteRewriteTunnelSmacRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_dmac_rewrite_req_ff.enq(req);
      end
    endcase
  endrule

  rule tunnel_src_rewrite_next_state if (tunnel_src_rewrite_rsp_ff.notEmpty);
    tunnel_src_rewrite_rsp_ff.deq;
    let _rsp = tunnel_src_rewrite_rsp_ff.first;
    case (_rsp) matches
      tagged TunnelSrcRewriteNopRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_dst_rewrite_req_ff.enq(req);
      end
      tagged TunnelSrcRewriteRewriteTunnelIpv4SrcRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_dst_rewrite_req_ff.enq(req);
      end
      tagged TunnelSrcRewriteRewriteTunnelIpv6SrcRspT {meta: .meta, pkt: .pkt}: begin
        MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
        tunnel_dst_rewrite_req_ff.enq(req);
      end
    endcase
  endrule

  rule vlan_decap_next_state if (vlan_decap_rsp_ff.notEmpty);
    vlan_decap_rsp_ff.deq;
    let _rsp = vlan_decap_rsp_ff.first;
    case (_rsp) matches
      tagged VlanDecapNopRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
        let multicast_metadata$replica = fromMaybe(?, meta.multicast_metadata$replica);
        let multicast_metadata$inner_replica = fromMaybe(?, meta.multicast_metadata$inner_replica);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( tunnel_metadata$tunnel_terminate == 'h1 )) begin
          if (( ( multicast_metadata$inner_replica == 'h1 ) || ( multicast_metadata$replica == 'h0 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_decap_process_outer_req_ff.enq(req);
          end
          else begin
            if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              rewrite_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              rewrite_multicast_req_ff.enq(req);
            end
          end
        end
        else begin
          if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            rewrite_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            rewrite_multicast_req_ff.enq(req);
          end
        end
      end
      tagged VlanDecapRemoveVlanSingleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
        let multicast_metadata$replica = fromMaybe(?, meta.multicast_metadata$replica);
        let multicast_metadata$inner_replica = fromMaybe(?, meta.multicast_metadata$inner_replica);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( tunnel_metadata$tunnel_terminate == 'h1 )) begin
          if (( ( multicast_metadata$inner_replica == 'h1 ) || ( multicast_metadata$replica == 'h0 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_decap_process_outer_req_ff.enq(req);
          end
          else begin
            if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              rewrite_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              rewrite_multicast_req_ff.enq(req);
            end
          end
        end
        else begin
          if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            rewrite_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            rewrite_multicast_req_ff.enq(req);
          end
        end
      end
      tagged VlanDecapRemoveVlanDoubleTaggedRspT {meta: .meta, pkt: .pkt}: begin
        let l3_metadata$nexthop_index = fromMaybe(?, meta.l3_metadata$nexthop_index);
        let multicast_metadata$replica = fromMaybe(?, meta.multicast_metadata$replica);
        let multicast_metadata$inner_replica = fromMaybe(?, meta.multicast_metadata$inner_replica);
        let tunnel_metadata$tunnel_terminate = fromMaybe(?, meta.tunnel_metadata$tunnel_terminate);
        let egress_metadata$routed = fromMaybe(?, meta.egress_metadata$routed);
        if (( tunnel_metadata$tunnel_terminate == 'h1 )) begin
          if (( ( multicast_metadata$inner_replica == 'h1 ) || ( multicast_metadata$replica == 'h0 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            tunnel_decap_process_outer_req_ff.enq(req);
          end
          else begin
            if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              rewrite_req_ff.enq(req);
            end
            else begin
              MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
              rewrite_multicast_req_ff.enq(req);
            end
          end
        end
        else begin
          if (( ( egress_metadata$routed == 'h0 ) || ( l3_metadata$nexthop_index != 'h0 ) )) begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            rewrite_req_ff.enq(req);
          end
          else begin
            MetadataRequest req = MetadataRequest {pkt: pkt, meta: meta};
            rewrite_multicast_req_ff.enq(req);
          end
        end
      end
    endcase
  endrule

  interface next = (interface Client#(MetadataRequest, MetadataResponse);
    interface request = toGet(next_req_ff);
    interface response = toPut(next_rsp_ff);
  endinterface);
endmodule
// Copyright (c) 2016 P4FPGA Project

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
