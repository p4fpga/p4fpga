typedef Bit#(36) ForwardReqSize;
typedef Bit#(50) ForwardRspSize;
typedef Bit#(36) Ipv4LpmReqSize;
typedef Bit#(43) Ipv4LpmRspSize;
typedef Bit#(9) SendFrameReqSize;
typedef Bit#(50) SendFrameRspSize;
