method forward_table_add_entry = prog.forward_table_add_entry;
method test_tbl_add_entry = prog.test_tbl_add_entry;
