import Ethernet::*;
typedef union tagged {
  struct {
    PacketInstance pkt;
  } Ipv4PacketReqT;
  struct {
    PacketInstance pkt;
  } Ipv6PacketReqT;
  struct {
    PacketInstance pkt;
  } L2PacketReqT;
  struct {
    PacketInstance pkt;
  } MimPacketReqT;
  struct {
    PacketInstance pkt;
  } MplsPacketReqT;
  struct {
    PacketInstance pkt;
  } NopReqT;
  struct {
    PacketInstance pkt;
    Bit#(8) runtime_egress_port_8;
  } SetEgressPortReqT;
} BBRequest deriving (Bits, Eq, FShow);
typedef union tagged {
  struct {
    PacketInstance pkt;
    Bit#(4) ing_metadata$packet_type;
  } Ipv4PacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ing_metadata$packet_type;
  } Ipv6PacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ing_metadata$packet_type;
  } L2PacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ing_metadata$packet_type;
  } MimPacketRspT;
  struct {
    PacketInstance pkt;
    Bit#(4) ing_metadata$packet_type;
  } MplsPacketRspT;
  struct {
    PacketInstance pkt;
  } NopRspT;
  struct {
    PacketInstance pkt;
    Bit#(8) ing_metadata$egress_port;
  } SetEgressPortRspT;
} BBResponse deriving (Bits, Eq, FShow);
