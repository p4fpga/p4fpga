//add more if need k>4

Vector#(4, G_Addr#(c, num_entries)) primes;

primes[0] = 997;
primes[1] = 79;
primes[2] = 267;
primes[3] = 533;
