import BUtils::*;
import BuildVector::*;
import CBus::*;
import ClientServer::*;
import ConfigReg::*;
import Connectable::*;
import DefaultValue::*;
import DbgDefs::*;
import FIFO::*;
import FIFOF::*;
import FShow::*;
import GetPut::*;
import List::*;
import MIMO::*;
import SpecialFIFOs::*;
import Vector::*;
import Ethernet::*;
import MatchTable::*;
import PacketBuffer::*;
import Pipe::*;
import PrintTrace::*;
import Register::*;
import StmtFSM::*;
import Stream::*;
import TxRx::*;
import TieOff::*;
import Utils::*;
import StructDefines::*;
import UnionDefines::*;

export BUtils::*;
export BuildVector::*;
export CBus::*;
export ClientServer::*;
export ConfigReg::*;
export Connectable::*;
export DefaultValue::*;
export DbgDefs::*;
export FIFO::*;
export FIFOF::*;
export FShow::*;
export GetPut::*;
export List::*;
export MIMO::*;
export SpecialFIFOs::*;
export Vector::*;
export Ethernet::*;
export MatchTable::*;
export PacketBuffer::*;
export Pipe::*;
export PrintTrace::*;
export Register::*;
export StmtFSM::*;
export Stream::*;
export TxRx::*;
export TieOff::*;
export Utils::*;
export StructDefines::*;
export UnionDefines::*;

