method forward_add_entry=prog.forward_add_entry;
// method ipv4_lpm_add_entry=ingress.ipv4_lpm_add_entry;
// method send_frame_add_entry=egress.send_frame_add_entry;
